module top(X0, X1, X2, X3, X4, X5, X6, X7, X8, X9, X10, out);
input [7:0] X0;
input [7:0] X1;
input [7:0] X2;
input [7:0] X3;
input [7:0] X4;
input [7:0] X5;
input [7:0] X6;
input [7:0] X7;
input [7:0] X8;
input [7:0] X9;
input [7:0] X10;
output [3:0] out;
assign out = 
   (X10 <= 84)?
     (X9 <= 38)?
       (X6 <= 39)?
         (X1 <= 80)?
           (X9 <= 22)?
            16
          :
             (X7 <= 106)?
               (X10 <= 32)?
                1
              :
                7
            :
               (X5 <= 63)?
                 (X5 <= 27)?
                   (X10 <= 55)?
                    10
                  :
                     (X10 <= 81)?
                       (X7 <= 137)?
                         (X4 <= 24)?
                          1
                        :
                          4
                      :
                        1
                    :
                      3
                :
                   (X1 <= 25)?
                    1
                  :
                     (X7 <= 107)?
                      2
                    :
                       (X6 <= 27)?
                         (X1 <= 55)?
                           (X6 <= 18)?
                            1
                          :
                            1
                        :
                          11
                      :
                         (X1 <= 50)?
                          3
                        :
                           (X3 <= 16)?
                             (X1 <= 53)?
                              1
                            :
                              2
                          :
                            3
              :
                 (X4 <= 27)?
                   (X5 <= 79)?
                    1
                  :
                    2
                :
                  3
        :
           (X0 <= 74)?
             (X1 <= 93)?
               (X2 <= 6)?
                3
              :
                 (X4 <= 31)?
                  4
                :
                  2
            :
               (X7 <= 90)?
                 (X4 <= 89)?
                  1
                :
                  1
              :
                 (X10 <= 69)?
                   (X6 <= 38)?
                    26
                  :
                    1
                :
                  1
          :
             (X6 <= 33)?
               (X9 <= 22)?
                 (X1 <= 103)?
                  7
                :
                   (X7 <= 100)?
                    1
                  :
                    5
              :
                 (X7 <= 136)?
                   (X7 <= 127)?
                     (X6 <= 22)?
                       (X7 <= 118)?
                        2
                      :
                        1
                    :
                      4
                  :
                    3
                :
                  12
            :
               (X2 <= 51)?
                3
              :
                 (X3 <= 22)?
                  2
                :
                   (X8 <= 96)?
                    1
                  :
                    1
      :
         (X10 <= 77)?
           (X5 <= 41)?
             (X3 <= 20)?
               (X8 <= 120)?
                1
              :
                1
            :
              13
          :
             (X3 <= 147)?
               (X6 <= 98)?
                 (X8 <= 161)?
                   (X2 <= 19)?
                    17
                  :
                     (X2 <= 73)?
                       (X8 <= 84)?
                        7
                      :
                         (X9 <= 34)?
                           (X8 <= 108)?
                             (X7 <= 125)?
                               (X1 <= 75)?
                                1
                              :
                                4
                            :
                              5
                          :
                             (X0 <= 56)?
                               (X0 <= 52)?
                                3
                              :
                                2
                            :
                              14
                        :
                          3
                    :
                       (X1 <= 19)?
                        1
                      :
                        20
                :
                  2
              :
                26
            :
              2
        :
           (X6 <= 75)?
            2
          :
             (X3 <= 123)?
              1
            :
              1
    :
       (X6 <= 69)?
         (X1 <= 53)?
           (X10 <= 53)?
             (X0 <= 138)?
               (X2 <= 137)?
                 (X8 <= 148)?
                   (X7 <= 118)?
                    2
                  :
                     (X4 <= 34)?
                       (X9 <= 39)?
                         (X8 <= 127)?
                          1
                        :
                          1
                      :
                        17
                    :
                       (X0 <= 78)?
                        2
                      :
                        3
                :
                  3
              :
                7
            :
              11
          :
             (X9 <= 71)?
               (X8 <= 75)?
                 (X7 <= 160)?
                  3
                :
                  2
              :
                 (X2 <= 105)?
                   (X0 <= 51)?
                     (X7 <= 91)?
                      1
                    :
                      5
                  :
                     (X4 <= 31)?
                       (X8 <= 99)?
                        1
                      :
                        7
                    :
                      2
                :
                   (X2 <= 124)?
                    8
                  :
                     (X5 <= 63)?
                       (X5 <= 25)?
                        2
                      :
                         (X10 <= 61)?
                          1
                        :
                          3
                    :
                      4
            :
               (X5 <= 20)?
                 (X4 <= 27)?
                  2
                :
                  3
              :
                 (X5 <= 49)?
                   (X4 <= 29)?
                     (X7 <= 150)?
                      1
                    :
                      3
                  :
                    2
                :
                  8
        :
           (X8 <= 161)?
             (X0 <= 121)?
               (X8 <= 112)?
                 (X10 <= 53)?
                   (X9 <= 192)?
                     (X2 <= 65)?
                      23
                    :
                       (X9 <= 48)?
                         (X0 <= 106)?
                          3
                        :
                          1
                      :
                         (X8 <= 42)?
                          1
                        :
                          12
                  :
                     (X1 <= 76)?
                      1
                    :
                      1
                :
                   (X9 <= 53)?
                     (X1 <= 95)?
                       (X10 <= 59)?
                        2
                      :
                        5
                    :
                      8
                  :
                    7
              :
                 (X1 <= 133)?
                   (X2 <= 81)?
                     (X10 <= 26)?
                      8
                    :
                       (X9 <= 72)?
                         (X8 <= 152)?
                           (X3 <= 36)?
                             (X10 <= 57)?
                               (X6 <= 38)?
                                 (X3 <= 18)?
                                   (X8 <= 135)?
                                     (X5 <= 59)?
                                       (X5 <= 34)?
                                         (X5 <= 9)?
                                          2
                                        :
                                           (X9 <= 53)?
                                            5
                                          :
                                            1
                                      :
                                         (X0 <= 62)?
                                          3
                                        :
                                          1
                                    :
                                      3
                                  :
                                    6
                                :
                                   (X1 <= 96)?
                                    12
                                  :
                                    4
                              :
                                10
                            :
                               (X6 <= 36)?
                                 (X8 <= 124)?
                                  5
                                :
                                   (X2 <= 3)?
                                    3
                                  :
                                     (X1 <= 75)?
                                      2
                                    :
                                       (X7 <= 125)?
                                         (X4 <= 69)?
                                          7
                                        :
                                          1
                                      :
                                         (X6 <= 25)?
                                          1
                                        :
                                          2
                              :
                                9
                          :
                            6
                        :
                           (X6 <= 21)?
                             (X7 <= 114)?
                              1
                            :
                               (X5 <= 41)?
                                2
                              :
                                1
                          :
                            7
                      :
                        8
                  :
                     (X5 <= 105)?
                      7
                    :
                      1
                :
                   (X3 <= 21)?
                    1
                  :
                    1
            :
               (X4 <= 54)?
                 (X8 <= 69)?
                   (X2 <= 140)?
                     (X3 <= 26)?
                       (X10 <= 72)?
                        2
                      :
                        1
                    :
                      2
                  :
                     (X9 <= 72)?
                      3
                    :
                      1
                :
                   (X5 <= 13)?
                    3
                  :
                     (X8 <= 87)?
                      8
                    :
                       (X9 <= 45)?
                        1
                      :
                         (X5 <= 96)?
                          6
                        :
                           (X7 <= 175)?
                            1
                          :
                            1
              :
                 (X5 <= 123)?
                  2
                :
                  1
          :
             (X5 <= 23)?
               (X7 <= 139)?
                 (X9 <= 45)?
                  2
                :
                  1
              :
                 (X9 <= 80)?
                  1
                :
                  2
            :
               (X3 <= 38)?
                16
              :
                1
      :
         (X9 <= 130)?
           (X3 <= 190)?
             (X1 <= 32)?
              1
            :
               (X9 <= 39)?
                 (X5 <= 85)?
                  2
                :
                  7
              :
                 (X3 <= 11)?
                  1
                :
                   (X6 <= 71)?
                     (X4 <= 26)?
                      1
                    :
                      3
                  :
                    48
          :
            2
        :
           (X10 <= 57)?
            2
          :
            4
  :
     (X9 <= 45)?
       (X1 <= 157)?
         (X1 <= 66)?
           (X8 <= 108)?
             (X7 <= 141)?
               (X3 <= 44)?
                 (X2 <= 106)?
                   (X6 <= 9)?
                    5
                  :
                     (X2 <= 92)?
                       (X10 <= 136)?
                        2
                      :
                        1
                    :
                      5
                :
                   (X10 <= 120)?
                     (X8 <= 97)?
                      1
                    :
                      1
                  :
                    9
              :
                5
            :
               (X4 <= 35)?
                3
              :
                3
          :
             (X7 <= 93)?
               (X7 <= 52)?
                 (X7 <= 48)?
                  3
                :
                  2
              :
                16
            :
               (X4 <= 25)?
                 (X10 <= 144)?
                  3
                :
                  2
              :
                 (X4 <= 29)?
                   (X8 <= 145)?
                    2
                  :
                    2
                :
                  5
        :
           (X5 <= 27)?
             (X3 <= 29)?
               (X7 <= 116)?
                 (X1 <= 72)?
                  1
                :
                   (X6 <= 5)?
                    3
                  :
                     (X1 <= 135)?
                       (X7 <= 38)?
                        1
                      :
                        7
                    :
                      2
              :
                 (X2 <= 27)?
                  2
                :
                  1
            :
              10
          :
             (X6 <= 12)?
               (X10 <= 126)?
                 (X7 <= 119)?
                  4
                :
                  1
              :
                4
            :
               (X9 <= 36)?
                 (X3 <= 46)?
                   (X5 <= 56)?
                    7
                  :
                     (X7 <= 76)?
                       (X6 <= 58)?
                        3
                      :
                        1
                    :
                       (X5 <= 106)?
                        4
                      :
                         (X10 <= 132)?
                          1
                        :
                          1
                :
                   (X1 <= 136)?
                    3
                  :
                    1
              :
                 (X5 <= 121)?
                   (X4 <= 18)?
                     (X7 <= 67)?
                      2
                    :
                      3
                  :
                     (X2 <= 87)?
                      24
                    :
                       (X7 <= 144)?
                        1
                      :
                        1
                :
                  2
      :
         (X3 <= 18)?
          2
        :
           (X9 <= 33)?
            3
          :
            3
    :
       (X10 <= 124)?
         (X1 <= 45)?
           (X6 <= 46)?
             (X8 <= 104)?
               (X0 <= 133)?
                 (X1 <= 39)?
                   (X8 <= 96)?
                    4
                  :
                    1
                :
                   (X2 <= 82)?
                    1
                  :
                    2
              :
                 (X1 <= 37)?
                  11
                :
                  1
            :
               (X6 <= 13)?
                 (X3 <= 22)?
                   (X9 <= 71)?
                    3
                  :
                    2
                :
                  3
              :
                 (X9 <= 62)?
                  6
                :
                   (X8 <= 131)?
                     (X8 <= 106)?
                       (X1 <= 35)?
                        1
                      :
                        2
                    :
                      5
                  :
                    5
          :
             (X0 <= 84)?
               (X4 <= 24)?
                 (X9 <= 86)?
                  2
                :
                  1
              :
                6
            :
               (X2 <= 143)?
                3
              :
                1
        :
           (X4 <= 35)?
             (X3 <= 25)?
               (X1 <= 91)?
                 (X8 <= 91)?
                   (X3 <= 24)?
                     (X6 <= 14)?
                      1
                    :
                      6
                  :
                    1
                :
                  28
              :
                 (X1 <= 94)?
                  3
                :
                  7
            :
               (X8 <= 117)?
                 (X9 <= 81)?
                  10
                :
                   (X9 <= 102)?
                    2
                  :
                    1
              :
                 (X7 <= 129)?
                   (X10 <= 96)?
                    3
                  :
                     (X1 <= 68)?
                      1
                    :
                      1
                :
                  5
          :
             (X0 <= 92)?
               (X3 <= 24)?
                3
              :
                1
            :
               (X6 <= 30)?
                7
              :
                 (X0 <= 127)?
                  2
                :
                  2
      :
         (X6 <= 12)?
           (X4 <= 32)?
             (X4 <= 24)?
               (X1 <= 46)?
                7
              :
                 (X9 <= 54)?
                  1
                :
                  4
            :
               (X6 <= 10)?
                 (X9 <= 51)?
                  1
                :
                  5
              :
                 (X1 <= 72)?
                  3
                :
                  1
          :
            10
        :
           (X9 <= 61)?
             (X8 <= 132)?
               (X5 <= 119)?
                15
              :
                1
            :
               (X4 <= 22)?
                 (X4 <= 15)?
                  2
                :
                   (X6 <= 25)?
                    1
                  :
                    2
              :
                 (X10 <= 140)?
                  1
                :
                  2
          :
             (X5 <= 63)?
               (X8 <= 100)?
                 (X7 <= 123)?
                  2
                :
                   (X10 <= 177)?
                    2
                  :
                    1
              :
                 (X1 <= 127)?
                   (X7 <= 133)?
                    20
                  :
                     (X8 <= 122)?
                      2
                    :
                      1
                :
                  1
            :
               (X8 <= 125)?
                 (X10 <= 215)?
                   (X4 <= 24)?
                    5
                  :
                     (X7 <= 123)?
                      5
                    :
                      4
                :
                  1
              :
                 (X6 <= 36)?
                   (X1 <= 74)?
                    2
                  :
                    1
                :
                  8
;
endmodule
