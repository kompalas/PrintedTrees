module top(X0, X1, X2, X3, X6, X7, X8, X9, X10, X11, X12, X13, X14, X15, X16, X17, X18, X19, out);
input [7:0] X0;
input [7:0] X1;
input [7:0] X2;
input [7:0] X3;
input [7:0] X6;
input [7:0] X7;
input [7:0] X8;
input [7:0] X9;
input [7:0] X10;
input [7:0] X11;
input [7:0] X12;
input [7:0] X13;
input [7:0] X14;
input [7:0] X15;
input [7:0] X16;
input [7:0] X17;
input [7:0] X18;
input [7:0] X19;
output [1:0] out;
assign out = 
   (X7[7:6] <= 3)?
     (X17[7:5] <= 3)?
       (X12[7:6] <= 1)?
         (X8[7:6] <= 2)?
          15
        :
          1
      :
         (X13[7:6] <= 1)?
          1
        :
          3
    :
       (X0[7:5] <= 5)?
         (X6[7:6] <= 0)?
           (X16[7:6] <= 0)?
            1
          :
             (X8[7:6] <= 0)?
               (X16[7:6] <= 1)?
                87
              :
                 (X0[7:6] <= 2)?
                   (X1[7:5] <= 0)?
                     (X17[7:6] <= 0)?
                      1
                    :
                      4
                  :
                    4
                :
                  32
            :
              535
        :
           (X2[7:6] <= 0)?
             (X10[7:6] <= 0)?
              31
            :
               (X14[7:6] <= 0)?
                1
              :
                1
          :
             (X1[7:6] <= 0)?
               (X13[7:5] <= 3)?
                1
              :
                3
            :
               (X19[7:6] <= 0)?
                6
              :
                 (X1[7:3] <= 4)?
                  2
                :
                  1
      :
         (X1[7:6] <= 0)?
           (X18[7:5] <= 3)?
             (X6[7:4] <= 1)?
               (X9[7:6] <= 1)?
                 (X2[7:6] <= 0)?
                  60
                :
                   (X2[7:5] <= 0)?
                    2
                  :
                    1
              :
                2
            :
              4
          :
             (X0[7:6] <= 1)?
               (X3[7:5] <= 0)?
                 (X18[7:5] <= 6)?
                  14
                :
                   (X11[7:6] <= 0)?
                    2
                  :
                    2
              :
                3
            :
               (X9[7:6] <= 2)?
                 (X13[7:6] <= 0)?
                   (X3[7:6] <= 0)?
                     (X15[7:6] <= 0)?
                      3
                    :
                       (X16[7:6] <= 0)?
                        1
                      :
                        1
                  :
                    16
                :
                   (X0[7:6] <= 1)?
                     (X7[7:6] <= 0)?
                       (X12[7:6] <= 4)?
                        4
                      :
                         (X1[7:6] <= 0)?
                          3
                        :
                          1
                    :
                      6
                  :
                     (X1[7:6] <= 0)?
                      6
                    :
                      1
              :
                4
        :
           (X3[7:6] <= 1)?
             (X9[7:4] <= 0)?
               (X19[7:6] <= 0)?
                2
              :
                33
            :
               (X10[7:5] <= 0)?
                1
              :
                3
          :
             (X15[7:6] <= 1)?
              144
            :
               (X12[7:6] <= 1)?
                5
              :
                1
  :
     (X9[7:6] <= 0)?
       (X17[7:5] <= 0)?
         (X13[7:6] <= 1)?
           (X14[7:6] <= 1)?
            45
          :
             (X6[7:4] <= 0)?
              1
            :
              1
        :
          2
      :
         (X7[7:6] <= 3)?
           (X19[7:6] <= 0)?
             (X12[7:5] <= 0)?
              5
            :
               (X3[7:5] <= 1)?
                 (X7[7:6] <= 1)?
                  2
                :
                  4
              :
                22
          :
             (X6[7:6] <= 0)?
              112
            :
               (X2[7:6] <= 0)?
                3
              :
                2
        :
           (X18[7:6] <= 1)?
            5
          :
            3
    :
       (X9[7:6] <= 1)?
         (X7[7:6] <= 1)?
           (X0[7:6] <= 1)?
             (X8[7:6] <= 0)?
               (X3[7:5] <= 1)?
                 (X1[7:5] <= 0)?
                   (X7[7:4] <= 13)?
                    26
                  :
                     (X9[7:6] <= 0)?
                      1
                    :
                      1
                :
                  2
              :
                 (X14[7:6] <= 0)?
                  4
                :
                  1
            :
               (X14[7:6] <= 0)?
                16
              :
                2
          :
             (X9[7:6] <= 0)?
               (X7[7:5] <= 3)?
                 (X9[7:6] <= 0)?
                   (X16[7:6] <= 0)?
                    37
                  :
                     (X1[7:5] <= 0)?
                      2
                    :
                      1
                :
                  1
              :
                 (X13[7:6] <= 0)?
                   (X2[7:6] <= 0)?
                    4
                  :
                    3
                :
                  4
            :
              82
        :
           (X3[7:5] <= 0)?
            8
          :
            2
      :
         (X3[7:6] <= 0)?
          24
        :
           (X8[7:6] <= 0)?
            1
          :
            2
;
endmodule
