module top(X0, X1, X2, X3, X4, X5, X6, X7, X8, X9, X10, out);
input [7:0] X0;
input [7:0] X1;
input [7:0] X2;
input [7:0] X3;
input [7:0] X4;
input [7:0] X5;
input [7:0] X6;
input [7:0] X7;
input [7:0] X8;
input [7:0] X9;
input [7:0] X10;
output [3:0] out;
assign out = 
   (X10[7:6] <= 1)?
     (X0[7:6] <= 0)?
       (X6[7:4] <= 3)?
         (X9[7:6] <= 0)?
           (X3[7:5] <= 0)?
             (X4[7:6] <= 0)?
               (X6[7:6] <= 0)?
                 (X2[7:6] <= 0)?
                   (X9[7:6] <= 0)?
                     (X0[7:6] <= 0)?
                       (X9[7:6] <= 0)?
                        13
                      :
                         (X0[7:5] <= 1)?
                           (X4[7:6] <= 0)?
                            1
                          :
                            5
                        :
                          2
                    :
                       (X10[7:6] <= 0)?
                        1
                      :
                        2
                  :
                    20
                :
                   (X1[7:6] <= 0)?
                    1
                  :
                     (X9[7:6] <= 0)?
                      1
                    :
                      4
              :
                3
            :
               (X4[7:4] <= 2)?
                 (X7[7:6] <= 0)?
                  20
                :
                   (X7[7:6] <= 1)?
                     (X0[7:6] <= 0)?
                      2
                    :
                      3
                  :
                    12
              :
                1
          :
             (X2[7:6] <= 0)?
              1
            :
              3
        :
           (X1[7:6] <= 0)?
             (X1[7:6] <= 0)?
              5
            :
               (X0[7:6] <= 0)?
                 (X1[7:6] <= 0)?
                   (X7[7:6] <= 0)?
                    3
                  :
                     (X6[7:5] <= 1)?
                       (X1[7:6] <= 0)?
                        7
                      :
                         (X10[7:5] <= 0)?
                          1
                        :
                          1
                    :
                      1
                :
                   (X0[7:5] <= 0)?
                    11
                  :
                     (X2[7:6] <= 0)?
                      8
                    :
                       (X6[7:6] <= 0)?
                         (X7[7:6] <= 1)?
                          7
                        :
                           (X7[7:6] <= 0)?
                             (X0[7:6] <= 0)?
                               (X4[7:6] <= 0)?
                                 (X8[7:6] <= 0)?
                                  11
                                :
                                   (X8[7:6] <= 0)?
                                    3
                                  :
                                     (X10[7:6] <= 0)?
                                      1
                                    :
                                       (X9[7:6] <= 0)?
                                        1
                                      :
                                        7
                              :
                                2
                            :
                              3
                          :
                             (X8[7:6] <= 0)?
                               (X7[7:4] <= 5)?
                                1
                              :
                                1
                            :
                              8
                      :
                         (X3[7:6] <= 0)?
                          14
                        :
                           (X0[7:6] <= 0)?
                             (X4[7:6] <= 0)?
                               (X4[7:6] <= 0)?
                                 (X1[7:6] <= 0)?
                                  1
                                :
                                  13
                              :
                                 (X1[7:6] <= 0)?
                                   (X2[7:6] <= 0)?
                                     (X1[7:5] <= 0)?
                                      2
                                    :
                                       (X0[7:6] <= 0)?
                                        3
                                      :
                                        1
                                  :
                                    4
                                :
                                  7
                            :
                              10
                          :
                             (X9[7:6] <= 0)?
                              1
                            :
                              8
              :
                 (X0[7:6] <= 0)?
                   (X9[7:6] <= 2)?
                     (X9[7:6] <= 0)?
                      18
                    :
                       (X0[7:6] <= 0)?
                        1
                      :
                        1
                  :
                     (X0[7:6] <= 1)?
                       (X9[7:4] <= 0)?
                        3
                      :
                         (X9[7:6] <= 0)?
                          7
                        :
                          1
                    :
                       (X7[7:5] <= 3)?
                        13
                      :
                         (X1[7:6] <= 0)?
                          1
                        :
                          2
                :
                   (X2[7:5] <= 3)?
                     (X0[7:6] <= 2)?
                      7
                    :
                      1
                  :
                    5
          :
             (X10[7:6] <= 0)?
              2
            :
               (X1[7:5] <= 0)?
                 (X0[7:6] <= 1)?
                   (X8[7:6] <= 0)?
                     (X5[7:6] <= 0)?
                       (X10[7:5] <= 0)?
                        2
                      :
                        1
                    :
                      8
                  :
                     (X7[7:6] <= 2)?
                       (X9[7:5] <= 0)?
                         (X5[7:6] <= 0)?
                          2
                        :
                          3
                      :
                         (X0[7:5] <= 0)?
                           (X4[7:6] <= 0)?
                             (X7[7:6] <= 0)?
                              6
                            :
                              1
                          :
                            2
                        :
                          13
                    :
                      13
                :
                   (X10[7:6] <= 0)?
                    3
                  :
                     (X2[7:6] <= 0)?
                      1
                    :
                      1
              :
                 (X9[7:5] <= 0)?
                  2
                :
                  2
      :
         (X4[7:6] <= 0)?
           (X6[7:6] <= 1)?
            2
          :
            3
        :
          45
    :
       (X9[7:6] <= 0)?
         (X1[7:5] <= 1)?
          5
        :
          1
      :
         (X5[7:6] <= 0)?
           (X9[7:6] <= 0)?
            13
          :
             (X0[7:4] <= 7)?
               (X9[7:5] <= 2)?
                1
              :
                3
            :
               (X7[7:6] <= 0)?
                1
              :
                2
        :
          2
  :
     (X9[7:6] <= 0)?
       (X10[7:6] <= 0)?
         (X6[7:5] <= 0)?
           (X1[7:6] <= 1)?
             (X3[7:6] <= 0)?
               (X8[7:6] <= 0)?
                 (X7[7:6] <= 0)?
                  5
                :
                   (X8[7:6] <= 0)?
                    1
                  :
                    2
              :
                 (X2[7:6] <= 0)?
                   (X8[7:6] <= 2)?
                    2
                  :
                     (X3[7:3] <= 0)?
                      1
                    :
                      1
                :
                  7
            :
               (X9[7:6] <= 0)?
                 (X1[7:6] <= 0)?
                   (X3[7:5] <= 0)?
                    5
                  :
                     (X0[7:5] <= 0)?
                       (X9[7:6] <= 1)?
                        4
                      :
                        2
                    :
                       (X0[7:5] <= 0)?
                        4
                      :
                         (X8[7:6] <= 0)?
                          6
                        :
                          1
                :
                   (X4[7:6] <= 0)?
                     (X6[7:6] <= 0)?
                      1
                    :
                       (X5[7:6] <= 1)?
                        15
                      :
                        1
                  :
                    1
              :
                 (X4[7:6] <= 0)?
                   (X10[7:6] <= 0)?
                    4
                  :
                     (X0[7:6] <= 2)?
                      1
                    :
                      1
                :
                   (X0[7:5] <= 0)?
                     (X6[7:6] <= 0)?
                      9
                    :
                      1
                  :
                    1
          :
             (X9[7:5] <= 0)?
               (X6[7:6] <= 0)?
                 (X1[7:5] <= 0)?
                   (X1[7:5] <= 1)?
                    1
                  :
                    3
                :
                  2
              :
                1
            :
               (X2[7:6] <= 0)?
                3
              :
                 (X7[7:6] <= 0)?
                  3
                :
                  1
        :
           (X9[7:6] <= 0)?
             (X10[7:6] <= 0)?
               (X3[7:6] <= 0)?
                 (X3[7:6] <= 0)?
                   (X4[7:5] <= 0)?
                    4
                  :
                    8
                :
                  25
              :
                 (X10[7:6] <= 0)?
                  2
                :
                  4
            :
               (X5[7:6] <= 0)?
                 (X2[7:4] <= 0)?
                   (X2[7:6] <= 0)?
                    1
                  :
                    2
                :
                  2
              :
                1
          :
             (X7[7:6] <= 0)?
               (X0[7:6] <= 0)?
                 (X1[7:6] <= 0)?
                   (X10[7:6] <= 0)?
                    1
                  :
                    4
                :
                   (X2[7:6] <= 0)?
                     (X5[7:6] <= 0)?
                       (X0[7:6] <= 2)?
                        19
                      :
                        1
                    :
                      2
                  :
                     (X2[7:6] <= 0)?
                       (X9[7:6] <= 0)?
                        8
                      :
                         (X6[7:6] <= 0)?
                          1
                        :
                          2
                    :
                       (X9[7:6] <= 0)?
                         (X5[7:6] <= 0)?
                           (X3[7:6] <= 0)?
                            4
                          :
                            3
                        :
                          9
                      :
                        2
              :
                 (X0[7:5] <= 1)?
                  1
                :
                  6
            :
              10
      :
         (X1[7:6] <= 0)?
           (X3[7:6] <= 0)?
             (X2[7:5] <= 4)?
               (X0[7:6] <= 0)?
                1
              :
                 (X4[7:6] <= 0)?
                  2
                :
                   (X6[7:5] <= 1)?
                     (X0[7:6] <= 0)?
                       (X0[7:6] <= 0)?
                         (X6[7:6] <= 0)?
                          1
                        :
                           (X6[7:6] <= 0)?
                            9
                          :
                             (X7[7:6] <= 0)?
                              1
                            :
                              1
                      :
                        3
                    :
                      8
                  :
                    20
            :
               (X8[7:5] <= 0)?
                1
              :
                1
          :
             (X2[7:6] <= 1)?
               (X7[7:6] <= 0)?
                1
              :
                2
            :
              5
        :
           (X7[7:5] <= 0)?
             (X8[7:6] <= 3)?
               (X2[7:6] <= 0)?
                 (X9[7:5] <= 0)?
                  3
                :
                  2
              :
                6
            :
              2
          :
             (X1[7:6] <= 1)?
               (X1[7:6] <= 0)?
                1
              :
                 (X4[7:6] <= 0)?
                  1
                :
                  7
            :
               (X1[7:6] <= 0)?
                1
              :
                1
    :
       (X10[7:3] <= 15)?
         (X1[7:6] <= 0)?
           (X6[7:6] <= 0)?
             (X8[7:6] <= 0)?
               (X0[7:6] <= 0)?
                 (X7[7:5] <= 2)?
                   (X10[7:6] <= 1)?
                    1
                  :
                    1
                :
                  2
              :
                 (X2[7:6] <= 2)?
                   (X3[7:6] <= 0)?
                     (X3[7:6] <= 0)?
                       (X6[7:5] <= 0)?
                         (X10[7:6] <= 0)?
                          7
                        :
                           (X1[7:4] <= 0)?
                            1
                          :
                            3
                      :
                         (X0[7:5] <= 0)?
                          3
                        :
                           (X7[7:5] <= 2)?
                             (X7[7:4] <= 5)?
                               (X2[7:6] <= 0)?
                                3
                              :
                                2
                            :
                              11
                          :
                            1
                    :
                       (X8[7:4] <= 2)?
                        1
                      :
                        1
                  :
                    6
                :
                  5
            :
               (X5[7:5] <= 0)?
                 (X9[7:6] <= 0)?
                   (X2[7:6] <= 0)?
                    3
                  :
                     (X2[7:6] <= 0)?
                       (X6[7:5] <= 0)?
                        1
                      :
                         (X6[7:5] <= 0)?
                           (X4[7:6] <= 0)?
                            2
                          :
                            1
                        :
                          2
                    :
                      5
                :
                   (X2[7:5] <= 1)?
                    8
                  :
                    1
              :
                 (X9[7:6] <= 0)?
                  10
                :
                   (X7[7:6] <= 1)?
                    5
                  :
                     (X7[7:5] <= 3)?
                       (X1[7:5] <= 0)?
                         (X10[7:6] <= 0)?
                          2
                        :
                          2
                      :
                        6
                    :
                      2
          :
             (X5[7:5] <= 0)?
               (X2[7:6] <= 1)?
                 (X8[7:5] <= 0)?
                  8
                :
                   (X2[7:6] <= 0)?
                    5
                  :
                    2
              :
                3
            :
               (X0[7:5] <= 2)?
                4
              :
                5
        :
           (X6[7:5] <= 0)?
             (X4[7:5] <= 0)?
               (X1[7:5] <= 0)?
                 (X1[7:5] <= 0)?
                   (X7[7:6] <= 1)?
                     (X7[7:5] <= 2)?
                       (X9[7:6] <= 1)?
                        8
                      :
                         (X7[7:5] <= 3)?
                          2
                        :
                          1
                    :
                      2
                  :
                     (X9[7:6] <= 0)?
                      1
                    :
                      12
                :
                   (X0[7:6] <= 0)?
                     (X8[7:4] <= 8)?
                      17
                    :
                      1
                  :
                     (X1[7:6] <= 0)?
                      3
                    :
                       (X8[7:6] <= 1)?
                        3
                      :
                         (X8[7:4] <= 4)?
                          20
                        :
                           (X2[7:5] <= 0)?
                            6
                          :
                            6
              :
                 (X1[7:6] <= 0)?
                  4
                :
                   (X10[7:6] <= 0)?
                     (X7[7:6] <= 0)?
                      5
                    :
                      3
                  :
                     (X1[7:6] <= 0)?
                      11
                    :
                      1
            :
               (X6[7:4] <= 0)?
                 (X2[7:6] <= 1)?
                   (X3[7:4] <= 0)?
                    2
                  :
                     (X3[7:6] <= 0)?
                       (X3[7:6] <= 0)?
                        4
                      :
                         (X5[7:4] <= 2)?
                          1
                        :
                          1
                    :
                      1
                :
                   (X2[7:6] <= 0)?
                     (X4[7:6] <= 0)?
                      12
                    :
                      1
                  :
                    2
              :
                6
          :
             (X9[7:6] <= 0)?
               (X2[7:6] <= 0)?
                 (X3[7:6] <= 0)?
                  1
                :
                   (X10[7:5] <= 0)?
                    1
                  :
                    1
              :
                15
            :
              4
      :
         (X10[7:6] <= 1)?
           (X9[7:6] <= 0)?
             (X6[7:5] <= 0)?
               (X3[7:6] <= 0)?
                1
              :
                6
            :
               (X3[7:6] <= 0)?
                 (X2[7:6] <= 0)?
                  1
                :
                  1
              :
                 (X0[7:6] <= 0)?
                   (X9[7:6] <= 0)?
                    14
                  :
                    1
                :
                  1
          :
             (X5[7:5] <= 1)?
               (X9[7:6] <= 0)?
                 (X0[7:6] <= 1)?
                  22
                :
                   (X3[7:6] <= 0)?
                    1
                  :
                    3
              :
                 (X5[7:6] <= 0)?
                   (X1[7:5] <= 0)?
                    1
                  :
                    5
                :
                  3
            :
               (X3[7:6] <= 0)?
                 (X10[7:5] <= 0)?
                  4
                :
                   (X2[7:6] <= 0)?
                    3
                  :
                     (X6[7:6] <= 0)?
                      4
                    :
                       (X6[7:6] <= 0)?
                        3
                      :
                         (X4[7:6] <= 0)?
                          2
                        :
                           (X8[7:5] <= 1)?
                             (X10[7:5] <= 0)?
                              2
                            :
                               (X4[7:6] <= 0)?
                                2
                              :
                                1
                          :
                            6
              :
                 (X10[7:5] <= 3)?
                  3
                :
                  1
        :
           (X6[7:6] <= 0)?
             (X4[7:6] <= 1)?
              2
            :
               (X9[7:6] <= 0)?
                3
              :
                2
          :
             (X5[7:6] <= 0)?
              2
            :
              3
;
endmodule
