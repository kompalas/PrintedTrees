
`timescale 1ns/1ps
module top_tb();
`define EOF 32'hFFFF_FFFF
`define NULL 0
localparam period = 0;
localparam halfperiod = period/2;

reg [7:0] X0_reg;
reg [7:0] X1_reg;
reg [7:0] X6_reg;
reg [7:0] X9_reg;
reg [7:0] X12_reg;
reg [7:0] X13_reg;
reg [7:0] X18_reg;
reg [7:0] X20_reg;
reg [7:0] X23_reg;
reg [7:0] X28_reg;
reg [7:0] X30_reg;
reg [7:0] X32_reg;
reg [7:0] X36_reg;
reg [7:0] X37_reg;
reg [7:0] X38_reg;
reg [7:0] X40_reg;
reg [7:0] X42_reg;
reg [7:0] X49_reg;
reg [7:0] X50_reg;
reg [7:0] X51_reg;
reg [7:0] X52_reg;
reg [7:0] X53_reg;
reg [7:0] X54_reg;
reg [7:0] X55_reg;
reg [7:0] X56_reg;
reg [7:0] X57_reg;
reg [7:0] X59_reg;
reg [7:0] X62_reg;
reg [7:0] X63_reg;
reg [7:0] X65_reg;
reg [7:0] X69_reg;
reg [7:0] X71_reg;
reg [7:0] X73_reg;
reg [7:0] X76_reg;
reg [7:0] X78_reg;
reg [7:0] X86_reg;
reg [7:0] X89_reg;
reg [7:0] X98_reg;
reg [7:0] X99_reg;
reg [7:0] X100_reg;
reg [7:0] X101_reg;
reg [7:0] X102_reg;
reg [7:0] X106_reg;
reg [7:0] X110_reg;
reg [7:0] X118_reg;
reg [7:0] X120_reg;
reg [7:0] X121_reg;
reg [7:0] X133_reg;
reg [7:0] X135_reg;
reg [7:0] X138_reg;
reg [7:0] X139_reg;
reg [7:0] X140_reg;
reg [7:0] X142_reg;
reg [7:0] X147_reg;
reg [7:0] X149_reg;
reg [7:0] X156_reg;
reg [7:0] X158_reg;
reg [7:0] X159_reg;
reg [7:0] X161_reg;
reg [7:0] X166_reg;
reg [7:0] X167_reg;
reg [7:0] X168_reg;
reg [7:0] X177_reg;
reg [7:0] X181_reg;
reg [7:0] X183_reg;
reg [7:0] X184_reg;
reg [7:0] X186_reg;
reg [7:0] X187_reg;
reg [7:0] X188_reg;
reg [7:0] X190_reg;
reg [7:0] X194_reg;
reg [7:0] X197_reg;
reg [7:0] X198_reg;
reg [7:0] X199_reg;
reg [7:0] X207_reg;
reg [7:0] X211_reg;
reg [7:0] X228_reg;
reg [7:0] X230_reg;
reg [7:0] X237_reg;
reg [7:0] X239_reg;
reg [7:0] X242_reg;
reg [7:0] X249_reg;
reg [7:0] X263_reg;
reg [7:0] X271_reg;
reg [7:0] X276_reg;
reg [7:0] X289_reg;
reg [7:0] X291_reg;
reg [7:0] X292_reg;
reg [7:0] X301_reg;
reg [7:0] X304_reg;
reg [7:0] X305_reg;
reg [7:0] X309_reg;
reg [7:0] X317_reg;
reg [7:0] X322_reg;
reg [7:0] X323_reg;
reg [7:0] X327_reg;
reg [7:0] X330_reg;
reg [7:0] X331_reg;
reg [7:0] X334_reg;
reg [7:0] X335_reg;
reg [7:0] X354_reg;
reg [7:0] X361_reg;
reg [7:0] X363_reg;
reg [7:0] X368_reg;
reg [7:0] X371_reg;
reg [7:0] X373_reg;
reg [7:0] X377_reg;
reg [7:0] X381_reg;
reg [7:0] X382_reg;
reg [7:0] X384_reg;
reg [7:0] X394_reg;
reg [7:0] X397_reg;
reg [7:0] X410_reg;
reg [7:0] X412_reg;
reg [7:0] X423_reg;
reg [7:0] X427_reg;
reg [7:0] X429_reg;
reg [7:0] X435_reg;
reg [7:0] X446_reg;
reg [7:0] X451_reg;
reg [7:0] X452_reg;
reg [7:0] X455_reg;
reg [7:0] X457_reg;
reg [7:0] X460_reg;
reg [7:0] X472_reg;
reg [7:0] X479_reg;
reg [7:0] X481_reg;
reg [7:0] X488_reg;
reg [7:0] X493_reg;
reg [7:0] X497_reg;
reg [7:0] X505_reg;
reg [7:0] X509_reg;
reg [7:0] X514_reg;
reg [7:0] X522_reg;
reg [7:0] X538_reg;
reg [7:0] X551_reg;
reg [7:0] X553_reg;
reg [7:0] X554_reg;
reg [7:0] X558_reg;
reg [7:0] X559_reg;
reg [7:0] X560_reg;
wire [7:0] X0;
wire [7:0] X1;
wire [7:0] X6;
wire [7:0] X9;
wire [7:0] X12;
wire [7:0] X13;
wire [7:0] X18;
wire [7:0] X20;
wire [7:0] X23;
wire [7:0] X28;
wire [7:0] X30;
wire [7:0] X32;
wire [7:0] X36;
wire [7:0] X37;
wire [7:0] X38;
wire [7:0] X40;
wire [7:0] X42;
wire [7:0] X49;
wire [7:0] X50;
wire [7:0] X51;
wire [7:0] X52;
wire [7:0] X53;
wire [7:0] X54;
wire [7:0] X55;
wire [7:0] X56;
wire [7:0] X57;
wire [7:0] X59;
wire [7:0] X62;
wire [7:0] X63;
wire [7:0] X65;
wire [7:0] X69;
wire [7:0] X71;
wire [7:0] X73;
wire [7:0] X76;
wire [7:0] X78;
wire [7:0] X86;
wire [7:0] X89;
wire [7:0] X98;
wire [7:0] X99;
wire [7:0] X100;
wire [7:0] X101;
wire [7:0] X102;
wire [7:0] X106;
wire [7:0] X110;
wire [7:0] X118;
wire [7:0] X120;
wire [7:0] X121;
wire [7:0] X133;
wire [7:0] X135;
wire [7:0] X138;
wire [7:0] X139;
wire [7:0] X140;
wire [7:0] X142;
wire [7:0] X147;
wire [7:0] X149;
wire [7:0] X156;
wire [7:0] X158;
wire [7:0] X159;
wire [7:0] X161;
wire [7:0] X166;
wire [7:0] X167;
wire [7:0] X168;
wire [7:0] X177;
wire [7:0] X181;
wire [7:0] X183;
wire [7:0] X184;
wire [7:0] X186;
wire [7:0] X187;
wire [7:0] X188;
wire [7:0] X190;
wire [7:0] X194;
wire [7:0] X197;
wire [7:0] X198;
wire [7:0] X199;
wire [7:0] X207;
wire [7:0] X211;
wire [7:0] X228;
wire [7:0] X230;
wire [7:0] X237;
wire [7:0] X239;
wire [7:0] X242;
wire [7:0] X249;
wire [7:0] X263;
wire [7:0] X271;
wire [7:0] X276;
wire [7:0] X289;
wire [7:0] X291;
wire [7:0] X292;
wire [7:0] X301;
wire [7:0] X304;
wire [7:0] X305;
wire [7:0] X309;
wire [7:0] X317;
wire [7:0] X322;
wire [7:0] X323;
wire [7:0] X327;
wire [7:0] X330;
wire [7:0] X331;
wire [7:0] X334;
wire [7:0] X335;
wire [7:0] X354;
wire [7:0] X361;
wire [7:0] X363;
wire [7:0] X368;
wire [7:0] X371;
wire [7:0] X373;
wire [7:0] X377;
wire [7:0] X381;
wire [7:0] X382;
wire [7:0] X384;
wire [7:0] X394;
wire [7:0] X397;
wire [7:0] X410;
wire [7:0] X412;
wire [7:0] X423;
wire [7:0] X427;
wire [7:0] X429;
wire [7:0] X435;
wire [7:0] X446;
wire [7:0] X451;
wire [7:0] X452;
wire [7:0] X455;
wire [7:0] X457;
wire [7:0] X460;
wire [7:0] X472;
wire [7:0] X479;
wire [7:0] X481;
wire [7:0] X488;
wire [7:0] X493;
wire [7:0] X497;
wire [7:0] X505;
wire [7:0] X509;
wire [7:0] X514;
wire [7:0] X522;
wire [7:0] X538;
wire [7:0] X551;
wire [7:0] X553;
wire [7:0] X554;
wire [7:0] X558;
wire [7:0] X559;
wire [7:0] X560;
wire [2:0] out;

integer fin, fout, r;

top DUT (X0, X1, X6, X9, X12, X13, X18, X20, X23, X28, X30, X32, X36, X37, X38, X40, X42, X49, X50, X51, X52, X53, X54, X55, X56, X57, X59, X62, X63, X65, X69, X71, X73, X76, X78, X86, X89, X98, X99, X100, X101, X102, X106, X110, X118, X120, X121, X133, X135, X138, X139, X140, X142, X147, X149, X156, X158, X159, X161, X166, X167, X168, X177, X181, X183, X184, X186, X187, X188, X190, X194, X197, X198, X199, X207, X211, X228, X230, X237, X239, X242, X249, X263, X271, X276, X289, X291, X292, X301, X304, X305, X309, X317, X322, X323, X327, X330, X331, X334, X335, X354, X361, X363, X368, X371, X373, X377, X381, X382, X384, X394, X397, X410, X412, X423, X427, X429, X435, X446, X451, X452, X455, X457, X460, X472, X479, X481, X488, X493, X497, X505, X509, X514, X522, X538, X551, X553, X554, X558, X559, X560, out);

//read inp
initial begin
    $display($time, " << Starting the Simulation >>");
    fin = $fopen("/home/balkon00/PrintedTrees/test/pareto/sim/inputs.txt", "r");
    if (fin == `NULL) begin
        $display($time, " file not found");
        $finish;
    end
    fout = $fopen("/home/balkon00/PrintedTrees/test/pareto/sim/output.txt", "w");
    forever begin
        r = $fscanf(fin,"%d\t%d\t%d\t%d\t%d\t%d\t%d\t%d\t%d\t%d\t%d\t%d\t%d\t%d\t%d\t%d\t%d\t%d\t%d\t%d\t%d\t%d\t%d\t%d\t%d\t%d\t%d\t%d\t%d\t%d\t%d\t%d\t%d\t%d\t%d\t%d\t%d\t%d\t%d\t%d\t%d\t%d\t%d\t%d\t%d\t%d\t%d\t%d\t%d\t%d\t%d\t%d\t%d\t%d\t%d\t%d\t%d\t%d\t%d\t%d\t%d\t%d\t%d\t%d\t%d\t%d\t%d\t%d\t%d\t%d\t%d\t%d\t%d\t%d\t%d\t%d\t%d\t%d\t%d\t%d\t%d\t%d\t%d\t%d\t%d\t%d\t%d\t%d\t%d\t%d\t%d\t%d\t%d\t%d\t%d\t%d\t%d\t%d\t%d\t%d\t%d\t%d\t%d\t%d\t%d\t%d\t%d\t%d\t%d\t%d\t%d\t%d\t%d\t%d\t%d\t%d\t%d\t%d\t%d\t%d\t%d\t%d\t%d\t%d\t%d\t%d\t%d\t%d\t%d\t%d\t%d\t%d\t%d\t%d\t%d\t%d\t%d\t%d\t%d\t%d\t%d\n", X0_reg, X1_reg, X6_reg, X9_reg, X12_reg, X13_reg, X18_reg, X20_reg, X23_reg, X28_reg, X30_reg, X32_reg, X36_reg, X37_reg, X38_reg, X40_reg, X42_reg, X49_reg, X50_reg, X51_reg, X52_reg, X53_reg, X54_reg, X55_reg, X56_reg, X57_reg, X59_reg, X62_reg, X63_reg, X65_reg, X69_reg, X71_reg, X73_reg, X76_reg, X78_reg, X86_reg, X89_reg, X98_reg, X99_reg, X100_reg, X101_reg, X102_reg, X106_reg, X110_reg, X118_reg, X120_reg, X121_reg, X133_reg, X135_reg, X138_reg, X139_reg, X140_reg, X142_reg, X147_reg, X149_reg, X156_reg, X158_reg, X159_reg, X161_reg, X166_reg, X167_reg, X168_reg, X177_reg, X181_reg, X183_reg, X184_reg, X186_reg, X187_reg, X188_reg, X190_reg, X194_reg, X197_reg, X198_reg, X199_reg, X207_reg, X211_reg, X228_reg, X230_reg, X237_reg, X239_reg, X242_reg, X249_reg, X263_reg, X271_reg, X276_reg, X289_reg, X291_reg, X292_reg, X301_reg, X304_reg, X305_reg, X309_reg, X317_reg, X322_reg, X323_reg, X327_reg, X330_reg, X331_reg, X334_reg, X335_reg, X354_reg, X361_reg, X363_reg, X368_reg, X371_reg, X373_reg, X377_reg, X381_reg, X382_reg, X384_reg, X394_reg, X397_reg, X410_reg, X412_reg, X423_reg, X427_reg, X429_reg, X435_reg, X446_reg, X451_reg, X452_reg, X455_reg, X457_reg, X460_reg, X472_reg, X479_reg, X481_reg, X488_reg, X493_reg, X497_reg, X505_reg, X509_reg, X514_reg, X522_reg, X538_reg, X551_reg, X553_reg, X554_reg, X558_reg, X559_reg, X560_reg);
        #period $fwrite(fout, "%d\n", out);
        if ($feof(fin)) begin
            $display($time, " << Finishing the Simulation >>");
            $fclose(fin);
            $fclose(fout);
            $finish;
        end
    end
end

assign X0 = X0_reg;
assign X1 = X1_reg;
assign X6 = X6_reg;
assign X9 = X9_reg;
assign X12 = X12_reg;
assign X13 = X13_reg;
assign X18 = X18_reg;
assign X20 = X20_reg;
assign X23 = X23_reg;
assign X28 = X28_reg;
assign X30 = X30_reg;
assign X32 = X32_reg;
assign X36 = X36_reg;
assign X37 = X37_reg;
assign X38 = X38_reg;
assign X40 = X40_reg;
assign X42 = X42_reg;
assign X49 = X49_reg;
assign X50 = X50_reg;
assign X51 = X51_reg;
assign X52 = X52_reg;
assign X53 = X53_reg;
assign X54 = X54_reg;
assign X55 = X55_reg;
assign X56 = X56_reg;
assign X57 = X57_reg;
assign X59 = X59_reg;
assign X62 = X62_reg;
assign X63 = X63_reg;
assign X65 = X65_reg;
assign X69 = X69_reg;
assign X71 = X71_reg;
assign X73 = X73_reg;
assign X76 = X76_reg;
assign X78 = X78_reg;
assign X86 = X86_reg;
assign X89 = X89_reg;
assign X98 = X98_reg;
assign X99 = X99_reg;
assign X100 = X100_reg;
assign X101 = X101_reg;
assign X102 = X102_reg;
assign X106 = X106_reg;
assign X110 = X110_reg;
assign X118 = X118_reg;
assign X120 = X120_reg;
assign X121 = X121_reg;
assign X133 = X133_reg;
assign X135 = X135_reg;
assign X138 = X138_reg;
assign X139 = X139_reg;
assign X140 = X140_reg;
assign X142 = X142_reg;
assign X147 = X147_reg;
assign X149 = X149_reg;
assign X156 = X156_reg;
assign X158 = X158_reg;
assign X159 = X159_reg;
assign X161 = X161_reg;
assign X166 = X166_reg;
assign X167 = X167_reg;
assign X168 = X168_reg;
assign X177 = X177_reg;
assign X181 = X181_reg;
assign X183 = X183_reg;
assign X184 = X184_reg;
assign X186 = X186_reg;
assign X187 = X187_reg;
assign X188 = X188_reg;
assign X190 = X190_reg;
assign X194 = X194_reg;
assign X197 = X197_reg;
assign X198 = X198_reg;
assign X199 = X199_reg;
assign X207 = X207_reg;
assign X211 = X211_reg;
assign X228 = X228_reg;
assign X230 = X230_reg;
assign X237 = X237_reg;
assign X239 = X239_reg;
assign X242 = X242_reg;
assign X249 = X249_reg;
assign X263 = X263_reg;
assign X271 = X271_reg;
assign X276 = X276_reg;
assign X289 = X289_reg;
assign X291 = X291_reg;
assign X292 = X292_reg;
assign X301 = X301_reg;
assign X304 = X304_reg;
assign X305 = X305_reg;
assign X309 = X309_reg;
assign X317 = X317_reg;
assign X322 = X322_reg;
assign X323 = X323_reg;
assign X327 = X327_reg;
assign X330 = X330_reg;
assign X331 = X331_reg;
assign X334 = X334_reg;
assign X335 = X335_reg;
assign X354 = X354_reg;
assign X361 = X361_reg;
assign X363 = X363_reg;
assign X368 = X368_reg;
assign X371 = X371_reg;
assign X373 = X373_reg;
assign X377 = X377_reg;
assign X381 = X381_reg;
assign X382 = X382_reg;
assign X384 = X384_reg;
assign X394 = X394_reg;
assign X397 = X397_reg;
assign X410 = X410_reg;
assign X412 = X412_reg;
assign X423 = X423_reg;
assign X427 = X427_reg;
assign X429 = X429_reg;
assign X435 = X435_reg;
assign X446 = X446_reg;
assign X451 = X451_reg;
assign X452 = X452_reg;
assign X455 = X455_reg;
assign X457 = X457_reg;
assign X460 = X460_reg;
assign X472 = X472_reg;
assign X479 = X479_reg;
assign X481 = X481_reg;
assign X488 = X488_reg;
assign X493 = X493_reg;
assign X497 = X497_reg;
assign X505 = X505_reg;
assign X509 = X509_reg;
assign X514 = X514_reg;
assign X522 = X522_reg;
assign X538 = X538_reg;
assign X551 = X551_reg;
assign X553 = X553_reg;
assign X554 = X554_reg;
assign X558 = X558_reg;
assign X559 = X559_reg;
assign X560 = X560_reg;

endmodule

