module top(X0, X1, X2, X3, X4, out);
input [7:0] X0;
input [7:0] X1;
input [7:0] X2;
input [7:0] X3;
input [7:0] X4;
output [0:0] out;
assign out = 
   (X0[7:1] <= 10)?
     (X2[7:4] <= 6)?
       (X1[7:4] <= 12)?
         (X3[7:2] <= 40)?
           (X4[7:3] <= 4)?
            1
          :
             (X1[7:5] <= 2)?
              42
            :
               (X1[7:3] <= 16)?
                 (X4[7:3] <= 15)?
                  17
                :
                   (X1[7:2] <= 30)?
                     (X1[7:5] <= 4)?
                       (X1[7:3] <= 8)?
                         (X1[7:3] <= 5)?
                           (X2[7:4] <= 3)?
                            3
                          :
                            2
                        :
                          17
                      :
                         (X0[7:4] <= 0)?
                          3
                        :
                           (X3[7:3] <= 4)?
                             (X1[7:2] <= 20)?
                               (X2[7:2] <= 11)?
                                3
                              :
                                4
                            :
                               (X2[7:3] <= 6)?
                                 (X1[7:3] <= 10)?
                                  2
                                :
                                  3
                              :
                                2
                          :
                            2
                    :
                       (X1[7:3] <= 13)?
                        40
                      :
                         (X1[7:5] <= 5)?
                           (X2[7:4] <= 3)?
                             (X1[7:5] <= 4)?
                              1
                            :
                              6
                          :
                            4
                        :
                          12
                  :
                     (X2[7:4] <= 0)?
                      2
                    :
                      1
              :
                22
        :
           (X1[7:5] <= 4)?
            5
          :
             (X3[7:3] <= 30)?
               (X2[7:4] <= 3)?
                1
              :
                 (X1[7:5] <= 8)?
                   (X1[7:4] <= 7)?
                    1
                  :
                    2
                :
                   (X1[7:4] <= 9)?
                     (X1[7:2] <= 35)?
                      1
                    :
                      1
                  :
                    2
            :
              1
      :
         (X1[7:5] <= 4)?
           (X1[7:4] <= 14)?
             (X2[7:6] <= 2)?
               (X4[7:3] <= 7)?
                1
              :
                 (X3[7:5] <= 4)?
                   (X3[7:4] <= 0)?
                     (X1[7:5] <= 8)?
                       (X1[7:5] <= 6)?
                        1
                      :
                         (X0[7:4] <= 2)?
                          1
                        :
                           (X1[7:3] <= 19)?
                            1
                          :
                            2
                    :
                      1
                  :
                    1
                :
                  1
            :
               (X3[7:3] <= 18)?
                5
              :
                1
          :
            2
        :
           (X4[7:2] <= 8)?
             (X1[7:3] <= 22)?
              1
            :
              1
          :
            9
    :
       (X1[7:3] <= 19)?
         (X1[7:3] <= 15)?
           (X1[7:5] <= 5)?
             (X1[7:4] <= 2)?
              2
            :
               (X1[7:4] <= 2)?
                1
              :
                 (X1[7:5] <= 3)?
                   (X1[7:5] <= 3)?
                     (X1[7:4] <= 5)?
                       (X3[7:4] <= 12)?
                        6
                      :
                        1
                    :
                       (X0[7:4] <= 0)?
                        1
                      :
                         (X3[7:4] <= 15)?
                           (X1[7:4] <= 10)?
                             (X3[7:4] <= 9)?
                               (X3[7:4] <= 4)?
                                 (X1[7:4] <= 7)?
                                  2
                                :
                                  2
                              :
                                 (X1[7:2] <= 27)?
                                  2
                                :
                                  1
                            :
                               (X1[7:6] <= 0)?
                                 (X4[7:3] <= 13)?
                                  1
                                :
                                  1
                              :
                                3
                          :
                            2
                        :
                          1
                  :
                     (X3[7:4] <= 14)?
                      6
                    :
                      1
                :
                   (X2[7:4] <= 11)?
                    1
                  :
                    2
          :
            6
        :
           (X1[7:3] <= 18)?
             (X1[7:5] <= 4)?
               (X4[7:3] <= 26)?
                 (X1[7:3] <= 15)?
                  1
                :
                   (X2[7:3] <= 28)?
                    1
                  :
                     (X3[7:4] <= 11)?
                      1
                    :
                      1
              :
                1
            :
               (X1[7:4] <= 9)?
                 (X3[7:4] <= 9)?
                  3
                :
                   (X1[7:3] <= 15)?
                    1
                  :
                     (X3[7:4] <= 15)?
                       (X2[7:5] <= 6)?
                        1
                      :
                        1
                    :
                      2
              :
                 (X3[7:3] <= 7)?
                  1
                :
                   (X4[7:4] <= 8)?
                    1
                  :
                     (X0[7:5] <= 2)?
                      1
                    :
                       (X3[7:3] <= 29)?
                         (X1[7:3] <= 18)?
                           (X3[7:3] <= 21)?
                            2
                          :
                             (X1[7:3] <= 18)?
                               (X2[7:5] <= 7)?
                                1
                              :
                                1
                            :
                              2
                        :
                           (X2[7:3] <= 28)?
                            2
                          :
                             (X1[7:2] <= 37)?
                               (X3[7:5] <= 5)?
                                1
                              :
                                1
                            :
                              1
                      :
                         (X1[7:4] <= 9)?
                          1
                        :
                          2
          :
            3
      :
         (X1[7:2] <= 46)?
           (X0[7:5] <= 0)?
            3
          :
             (X1[7:3] <= 23)?
               (X1[7:2] <= 42)?
                 (X1[7:4] <= 9)?
                   (X3[7:3] <= 12)?
                    1
                  :
                     (X1[7:4] <= 9)?
                       (X3[7:4] <= 15)?
                        2
                      :
                        1
                    :
                       (X3[7:2] <= 59)?
                        2
                      :
                        1
                :
                  1
              :
                6
            :
               (X4[7:4] <= 8)?
                1
              :
                 (X3[7:4] <= 4)?
                  1
                :
                   (X3[7:5] <= 2)?
                    1
                  :
                     (X2[7:4] <= 15)?
                      1
                    :
                       (X3[7:4] <= 9)?
                         (X1[7:3] <= 23)?
                          1
                        :
                          1
                      :
                        1
        :
          4
  :
     (X4[7:3] <= 27)?
       (X3[7:4] <= 2)?
         (X0[7:3] <= 3)?
           (X2[7:3] <= 18)?
            5
          :
             (X4[7:4] <= 2)?
              1
            :
              1
        :
          2
      :
         (X1[7:4] <= 1)?
           (X2[7:4] <= 11)?
            1
          :
            1
        :
           (X4 <= 127)?
             (X2[7:4] <= 7)?
              1
            :
               (X1[7:4] <= 10)?
                 (X1[7:4] <= 9)?
                  3
                :
                  1
              :
                4
          :
             (X1[7:4] <= 16)?
               (X1[7:4] <= 10)?
                 (X1[7:4] <= 10)?
                   (X1[7:3] <= 10)?
                     (X1[7:5] <= 2)?
                      5
                    :
                       (X3[7:4] <= 12)?
                        1
                      :
                        1
                  :
                    27
                :
                   (X1[7:5] <= 4)?
                     (X2[7:2] <= 53)?
                      1
                    :
                       (X1[7:4] <= 7)?
                         (X3[7:2] <= 46)?
                          1
                        :
                          1
                      :
                         (X3[7:3] <= 20)?
                          1
                        :
                          3
                  :
                     (X1[7:4] <= 11)?
                      10
                    :
                       (X1[7:3] <= 15)?
                         (X2[7:3] <= 21)?
                          1
                        :
                          1
                      :
                         (X3[7:3] <= 13)?
                           (X1[7:3] <= 20)?
                            1
                          :
                            3
                        :
                           (X1[7:4] <= 8)?
                            19
                          :
                             (X3[7:6] <= 2)?
                              15
                            :
                               (X1[7:3] <= 22)?
                                 (X1[7:5] <= 5)?
                                   (X1[7:3] <= 18)?
                                     (X3[7:1] <= 109)?
                                      1
                                    :
                                      2
                                  :
                                     (X1[7:4] <= 7)?
                                      6
                                    :
                                       (X3[7:3] <= 27)?
                                         (X1[7:1] <= 77)?
                                          2
                                        :
                                          6
                                      :
                                         (X1[7:3] <= 19)?
                                          3
                                        :
                                          1
                                :
                                   (X1[7:6] <= 4)?
                                    18
                                  :
                                     (X3[7:4] <= 14)?
                                      4
                                    :
                                      2
                              :
                                 (X2[7:3] <= 23)?
                                  1
                                :
                                  1
              :
                41
            :
               (X1[7:5] <= 7)?
                 (X2[7:6] <= 1)?
                  2
                :
                   (X1[7:5] <= 6)?
                     (X3[7:5] <= 8)?
                      3
                    :
                      1
                  :
                    1
              :
                6
    :
       (X1[7:4] <= 6)?
        1
      :
         (X3[7:5] <= 4)?
          1
        :
           (X1[7:4] <= 9)?
            1
          :
             (X1[7:6] <= 0)?
              1
            :
              1
;
endmodule
