module top(X0, X1, X2, X3, X4, X5, X6, X7, X8, X9, X10, X11, X12, X13, X14, X15, out);
input [7:0] X0;
input [7:0] X1;
input [7:0] X2;
input [7:0] X3;
input [7:0] X4;
input [7:0] X5;
input [7:0] X6;
input [7:0] X7;
input [7:0] X8;
input [7:0] X9;
input [7:0] X10;
input [7:0] X11;
input [7:0] X12;
input [7:0] X13;
input [7:0] X14;
input [7:0] X15;
output [3:0] out;
assign out = 
   (X15[7:3] <= 8)?
     (X4[7:5] <= 3)?
       (X9[7:5] <= 2)?
         (X14[7:3] <= 15)?
          349
        :
           (X13[7:5] <= 0)?
             (X12[7:6] <= 2)?
              19
            :
              21
          :
             (X9[7:4] <= 0)?
              1
            :
              28
      :
         (X5[7:5] <= 4)?
           (X7[7:5] <= 6)?
             (X15[7:6] <= 0)?
               (X5[7:3] <= 3)?
                2
              :
                 (X9[7:6] <= 1)?
                  682
                :
                   (X11[7:6] <= 0)?
                    1
                  :
                    8
            :
               (X5[7:5] <= 3)?
                17
              :
                2
          :
             (X10[7:6] <= 3)?
               (X0[7:5] <= 6)?
                 (X13[7:4] <= 0)?
                   (X12[7:5] <= 2)?
                    1
                  :
                    1
                :
                  21
              :
                 (X13[7:5] <= 2)?
                  4
                :
                  1
            :
              38
        :
           (X9[7:5] <= 6)?
             (X14[7:4] <= 1)?
               (X6[7:5] <= 4)?
                 (X10[7:5] <= 2)?
                   (X7[7:5] <= 4)?
                    1
                  :
                    4
                :
                   (X2[7:4] <= 6)?
                     (X0[7:6] <= 0)?
                      2
                    :
                       (X5[7:5] <= 3)?
                        1
                      :
                        1
                  :
                     (X1[7:3] <= 21)?
                      1
                    :
                      91
              :
                 (X9[7:5] <= 1)?
                   (X0[7:4] <= 14)?
                    1
                  :
                    7
                :
                  33
            :
               (X10[7:5] <= 3)?
                 (X12[7:6] <= 0)?
                  19
                :
                   (X7[7:5] <= 5)?
                    6
                  :
                    1
              :
                 (X9[7:5] <= 5)?
                   (X13[7:4] <= 1)?
                     (X8[7:6] <= 0)?
                       (X6[7:5] <= 0)?
                        1
                      :
                        1
                    :
                      3
                  :
                    56
                :
                   (X5[7:5] <= 5)?
                    2
                  :
                    7
          :
             (X0[7:5] <= 0)?
               (X7[7:5] <= 6)?
                 (X11[7:6] <= 0)?
                   (X3[7:5] <= 8)?
                    1
                  :
                    3
                :
                  3
              :
                 (X1[7:3] <= 17)?
                  3
                :
                  24
            :
               (X1[7:4] <= 12)?
                207
              :
                 (X7[7:4] <= 10)?
                   (X13[7:4] <= 2)?
                    1
                  :
                    5
                :
                   (X5[7:6] <= 4)?
                    29
                  :
                    2
    :
       (X14[7:5] <= 2)?
         (X3[7:4] <= 15)?
           (X10[7:3] <= 23)?
             (X7[7:5] <= 4)?
               (X9[7:3] <= 10)?
                13
              :
                 (X5[7:6] <= 2)?
                  11
                :
                  1
            :
               (X0[7:5] <= 2)?
                 (X8[7:5] <= 0)?
                   (X13[7:5] <= 2)?
                     (X12[7:3] <= 6)?
                      1
                    :
                       (X1[7:3] <= 12)?
                        1
                      :
                        1
                  :
                    6
                :
                   (X3[7:3] <= 27)?
                     (X2[7:6] <= 0)?
                       (X3[7:4] <= 12)?
                         (X4[7:6] <= 0)?
                          5
                        :
                          1
                      :
                        2
                    :
                       (X13[7:2] <= 28)?
                        211
                      :
                        1
                  :
                     (X2[7:3] <= 7)?
                      9
                    :
                      4
              :
                 (X10[7:6] <= 2)?
                   (X3[7:5] <= 5)?
                     (X5[7:6] <= 3)?
                      2
                    :
                       (X5[7:5] <= 4)?
                        1
                      :
                        1
                  :
                    43
                :
                   (X0[7:4] <= 4)?
                     (X9[7:6] <= 0)?
                      5
                    :
                       (X3[7:5] <= 3)?
                         (X2[7:4] <= 3)?
                          1
                        :
                          1
                      :
                        3
                  :
                     (X7[7:6] <= 1)?
                      1
                    :
                      29
          :
             (X1[7:3] <= 18)?
               (X6[7:6] <= 1)?
                 (X13[7:6] <= 1)?
                  6
                :
                  4
              :
                11
            :
               (X9[7:5] <= 2)?
                 (X0[7:5] <= 3)?
                  2
                :
                  3
              :
                 (X0[7:5] <= 0)?
                   (X3[7:5] <= 5)?
                    10
                  :
                     (X2[7:5] <= 3)?
                      3
                    :
                       (X2[7:6] <= 3)?
                        2
                      :
                        1
                :
                   (X9[7:6] <= 1)?
                     (X0[7:4] <= 10)?
                      2
                    :
                      5
                  :
                    163
        :
           (X7[7:3] <= 25)?
             (X2[7:3] <= 29)?
               (X4[7:4] <= 9)?
                 (X9[7:5] <= 2)?
                   (X0[7:5] <= 2)?
                    2
                  :
                    7
                :
                   (X6[7:6] <= 3)?
                     (X2[7:4] <= 7)?
                      6
                    :
                       (X14[7:5] <= 3)?
                         (X1[7:4] <= 13)?
                          1
                        :
                           (X10[7:4] <= 1)?
                            1
                          :
                            23
                      :
                        2
                  :
                    9
              :
                 (X12[7:5] <= 3)?
                   (X15[7:3] <= 4)?
                    6
                  :
                     (X13[7:6] <= 0)?
                      1
                    :
                      3
                :
                   (X9[7:3] <= 6)?
                     (X15[7:6] <= 1)?
                      3
                    :
                       (X14[7:5] <= 1)?
                        1
                      :
                        2
                  :
                     (X3[7:2] <= 59)?
                       (X0[7:5] <= 7)?
                         (X6[7:6] <= 4)?
                           (X6[7:3] <= 12)?
                            1
                          :
                            16
                        :
                           (X1[7:5] <= 4)?
                            2
                          :
                            3
                      :
                         (X1[7:6] <= 4)?
                          1
                        :
                          3
                    :
                       (X5[7:5] <= 4)?
                        1
                      :
                         (X13[7:5] <= 2)?
                           (X2[7:6] <= 2)?
                            643
                          :
                             (X13[7:4] <= 3)?
                              16
                            :
                              1
                        :
                           (X10[7:4] <= 11)?
                            1
                          :
                            1
            :
               (X5[7:6] <= 1)?
                 (X13[7:5] <= 0)?
                   (X4[7:5] <= 4)?
                     (X2[7:3] <= 31)?
                      2
                    :
                      9
                  :
                     (X10[7:5] <= 2)?
                      2
                    :
                      23
                :
                   (X9[7:3] <= 11)?
                     (X9[7:4] <= 4)?
                      11
                    :
                      1
                  :
                    20
              :
                 (X1[7:3] <= 23)?
                  8
                :
                   (X6[7:4] <= 10)?
                     (X11[7:5] <= 4)?
                      64
                    :
                      1
                  :
                     (X15[7:6] <= 0)?
                       (X11[7:5] <= 3)?
                        1
                      :
                        2
                    :
                      2
          :
             (X5[7:4] <= 14)?
              92
            :
               (X2[7:5] <= 4)?
                 (X11[7:4] <= 5)?
                   (X10[7:5] <= 5)?
                    2
                  :
                    25
                :
                   (X2[7:6] <= 2)?
                    55
                  :
                     (X1[7:3] <= 30)?
                       (X1[7:4] <= 13)?
                        1
                      :
                         (X14[7:3] <= 4)?
                          1
                        :
                          1
                    :
                      4
              :
                 (X13[7:4] <= 0)?
                   (X11[7:4] <= 0)?
                    1
                  :
                    76
                :
                   (X11[7:3] <= 14)?
                    2
                  :
                    1
      :
         (X3[7:4] <= 13)?
           (X6[7:4] <= 6)?
             (X9[7:5] <= 0)?
               (X14[7:5] <= 8)?
                1
              :
                1
            :
              38
          :
             (X8[7:5] <= 3)?
               (X8[7:6] <= 2)?
                6
              :
                1
            :
               (X1[7:3] <= 30)?
                 (X10[7:5] <= 0)?
                   (X6[7:6] <= 0)?
                    12
                  :
                    4
                :
                   (X13[7:4] <= 6)?
                    257
                  :
                    1
              :
                 (X14[7:6] <= 2)?
                  3
                :
                  1
        :
           (X8[7:3] <= 7)?
             (X9[7:3] <= 3)?
               (X8[7:3] <= 1)?
                 (X4[7:5] <= 3)?
                   (X0[7:5] <= 1)?
                    15
                  :
                     (X5[7:3] <= 22)?
                      4
                    :
                      4
                :
                  105
              :
                 (X4[7:5] <= 5)?
                   (X8[7:5] <= 2)?
                     (X7[7:3] <= 8)?
                       (X12[7:6] <= 2)?
                        1
                      :
                        2
                    :
                       (X7[7:3] <= 14)?
                        7
                      :
                        1
                  :
                    15
                :
                   (X1[7:4] <= 11)?
                    26
                  :
                     (X6[7:6] <= 2)?
                      3
                    :
                      1
            :
               (X9[7:6] <= 2)?
                 (X5[7:3] <= 29)?
                  335
                :
                   (X2[7:6] <= 0)?
                    56
                  :
                     (X4[7:5] <= 5)?
                      3
                    :
                      25
              :
                 (X10[7:4] <= 7)?
                  2
                :
                  1
          :
             (X15[7:4] <= 3)?
               (X6[7:5] <= 3)?
                 (X2[7:4] <= 3)?
                  18
                :
                   (X13[7:4] <= 0)?
                    80
                  :
                     (X2[7:3] <= 13)?
                      3
                    :
                      7
              :
                 (X8[7:4] <= 11)?
                   (X2[7:5] <= 4)?
                    108
                  :
                     (X4[7:4] <= 12)?
                       (X5[7:4] <= 10)?
                        2
                      :
                        16
                    :
                       (X8[7:6] <= 2)?
                         (X0[7:3] <= 0)?
                           (X2[7:6] <= 2)?
                            2
                          :
                            1
                        :
                          46
                      :
                         (X2[7:5] <= 4)?
                          2
                        :
                          3
                :
                   (X2[7:5] <= 3)?
                     (X14[7:4] <= 10)?
                       (X1[7:5] <= 4)?
                        1
                      :
                        8
                    :
                       (X7[7:4] <= 11)?
                        1
                      :
                        4
                  :
                    15
            :
               (X0[7:3] <= 4)?
                27
              :
                1
  :
     (X13[7:4] <= 12)?
       (X0[7:6] <= 1)?
         (X14[7:3] <= 16)?
           (X1[7:6] <= 2)?
             (X8[7:4] <= 11)?
               (X12[7:4] <= 14)?
                34
              :
                 (X5[7:6] <= 3)?
                  1
                :
                  2
            :
              5
          :
             (X3[7:5] <= 5)?
               (X4[7:6] <= 1)?
                2
              :
                8
            :
               (X9[7:4] <= 5)?
                 (X15[7:5] <= 3)?
                  59
                :
                   (X11[7:4] <= 0)?
                    1
                  :
                    1
              :
                2
        :
           (X8[7:6] <= 0)?
             (X0[7:2] <= 5)?
              1
            :
              13
          :
             (X1[7:4] <= 11)?
               (X15[7:5] <= 3)?
                 (X2[7:4] <= 7)?
                  6
                :
                  1
              :
                2
            :
              563
      :
         (X6[7:3] <= 10)?
           (X14[7:3] <= 17)?
             (X9[7:4] <= 6)?
               (X15[7:5] <= 6)?
                324
              :
                1
            :
               (X13[7:4] <= 1)?
                 (X11[7:4] <= 3)?
                  4
                :
                  2
              :
                 (X15[7:3] <= 6)?
                  1
                :
                  12
          :
             (X12[7:4] <= 9)?
              17
            :
              29
        :
           (X15[7:3] <= 11)?
             (X7[7:5] <= 5)?
               (X10[7:6] <= 1)?
                 (X2[7:5] <= 3)?
                  1
                :
                  4
              :
                 (X0[7:3] <= 16)?
                  2
                :
                  3
            :
               (X11[7:4] <= 0)?
                 (X3[7:6] <= 4)?
                   (X4[7:4] <= 4)?
                    1
                  :
                    3
                :
                  4
              :
                6
          :
             (X15[7:3] <= 16)?
               (X7[7:5] <= 3)?
                3
              :
                17
            :
              177
    :
       (X8[7:4] <= 8)?
         (X14[7:5] <= 6)?
           (X12[7:6] <= 0)?
            9
          :
             (X11[7:5] <= 1)?
               (X12[7:4] <= 15)?
                16
              :
                12
            :
               (X1[7:4] <= 6)?
                1
              :
                331
        :
           (X13[7:4] <= 13)?
             (X6[7:5] <= 0)?
              4
            :
               (X11[7:5] <= 4)?
                 (X5[7:5] <= 4)?
                   (X9[7:5] <= 0)?
                    1
                  :
                    1
                :
                  40
              :
                 (X5[7:4] <= 6)?
                  3
                :
                  1
          :
             (X12[7:5] <= 6)?
               (X5[7:3] <= 17)?
                377
              :
                 (X12[7:4] <= 7)?
                  47
                :
                  1
            :
              1
      :
         (X7[7:5] <= 3)?
           (X2[7:5] <= 4)?
             (X6[7:4] <= 15)?
               (X4[7:4] <= 7)?
                716
              :
                 (X3[7:4] <= 6)?
                  1
                :
                  1
            :
               (X15[7:6] <= 2)?
                11
              :
                4
          :
             (X11[7:6] <= 0)?
               (X6[7:5] <= 0)?
                1
              :
                1
            :
              11
        :
           (X9[7:5] <= 2)?
             (X12[7:4] <= 2)?
              1
            :
              31
          :
             (X5[7:6] <= 1)?
               (X6[7:6] <= 2)?
                2
              :
                24
            :
              16
;
endmodule
