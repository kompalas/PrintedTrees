module top(X0, X1, X2, X3, X4, X5, X6, X7, X8, X9, X10, out);
input [7:0] X0;
input [7:0] X1;
input [7:0] X2;
input [7:0] X3;
input [7:0] X4;
input [7:0] X5;
input [7:0] X6;
input [7:0] X7;
input [7:0] X8;
input [7:0] X9;
input [7:0] X10;
output [3:0] out;
assign out = 
   (X10[7:3] <= 11)?
     (X0[7:1] <= 70)?
       (X6[7:4] <= 4)?
         (X9[7:3] <= 4)?
           (X3[7:4] <= 7)?
             (X4[7:2] <= 8)?
               (X6[7:4] <= 7)?
                 (X2[7:3] <= 10)?
                   (X9[7:3] <= 4)?
                     (X0[7:3] <= 9)?
                       (X9[7:4] <= 3)?
                        13
                      :
                         (X0[7:4] <= 6)?
                           (X4[7:3] <= 1)?
                            1
                          :
                            5
                        :
                          2
                    :
                       (X10[7:3] <= 7)?
                        1
                      :
                        2
                  :
                    20
                :
                   (X1[7:3] <= 3)?
                    1
                  :
                     (X9[7:3] <= 3)?
                      1
                    :
                      4
              :
                3
            :
               (X4[7:3] <= 9)?
                 (X7[7:3] <= 18)?
                  20
                :
                   (X7[7:5] <= 4)?
                     (X0[7:4] <= 6)?
                      2
                    :
                      3
                  :
                    12
              :
                1
          :
             (X2[7:3] <= 7)?
              1
            :
              3
        :
           (X1[7:1] <= 46)?
             (X1[7:2] <= 4)?
              5
            :
               (X0[7:5] <= 3)?
                 (X1[7:3] <= 5)?
                   (X7[7:3] <= 15)?
                    3
                  :
                     (X6[7:4] <= 5)?
                       (X1[7:3] <= 6)?
                        7
                      :
                         (X10[7:5] <= 0)?
                          1
                        :
                          1
                    :
                      1
                :
                   (X0[7:2] <= 11)?
                    11
                  :
                     (X2[7:4] <= 0)?
                      8
                    :
                       (X6[7:3] <= 5)?
                         (X7[7:3] <= 14)?
                          7
                        :
                           (X7[7:1] <= 72)?
                             (X0[7:1] <= 37)?
                               (X4[7:3] <= 8)?
                                 (X8[7:2] <= 28)?
                                  11
                                :
                                   (X8[7:2] <= 34)?
                                    3
                                  :
                                     (X10[7:3] <= 5)?
                                      1
                                    :
                                       (X9[7:2] <= 13)?
                                        1
                                      :
                                        7
                              :
                                2
                            :
                              3
                          :
                             (X8[7:2] <= 26)?
                               (X7[7:3] <= 19)?
                                1
                              :
                                1
                            :
                              8
                      :
                         (X3[7:6] <= 0)?
                          14
                        :
                           (X0[7:4] <= 6)?
                             (X4[7:2] <= 4)?
                               (X4[7:4] <= 1)?
                                 (X1[7:3] <= 6)?
                                  1
                                :
                                  13
                              :
                                 (X1[7:2] <= 20)?
                                   (X2[7:4] <= 7)?
                                     (X1[7:4] <= 2)?
                                      2
                                    :
                                       (X0[7:2] <= 20)?
                                        3
                                      :
                                        1
                                  :
                                    4
                                :
                                  7
                            :
                              10
                          :
                             (X9[7:4] <= 3)?
                              1
                            :
                              8
              :
                 (X0[7:5] <= 4)?
                   (X9[7:4] <= 3)?
                     (X9[7:3] <= 6)?
                      18
                    :
                       (X0[7:3] <= 17)?
                        1
                      :
                        1
                  :
                     (X0[7:3] <= 12)?
                       (X9[7:2] <= 13)?
                        3
                      :
                         (X9[7:1] <= 81)?
                          7
                        :
                          1
                    :
                       (X7[7:2] <= 54)?
                        13
                      :
                         (X1[7:3] <= 8)?
                          1
                        :
                          2
                :
                   (X2[7:5] <= 5)?
                     (X0[7:1] <= 67)?
                      7
                    :
                      1
                  :
                    5
          :
             (X10[7:2] <= 7)?
              2
            :
               (X1[7:3] <= 16)?
                 (X0[7:2] <= 25)?
                   (X8[7:4] <= 6)?
                     (X5[7:2] <= 10)?
                       (X10[7:5] <= 1)?
                        2
                      :
                        1
                    :
                      8
                  :
                     (X7[7:5] <= 4)?
                       (X9[7:2] <= 8)?
                         (X5[7:2] <= 7)?
                          2
                        :
                          3
                      :
                         (X0[7:2] <= 14)?
                           (X4[7:4] <= 1)?
                             (X7[7:5] <= 3)?
                              6
                            :
                              1
                          :
                            2
                        :
                          13
                    :
                      13
                :
                   (X10[7:5] <= 1)?
                    3
                  :
                     (X2[7:2] <= 6)?
                      1
                    :
                      1
              :
                 (X9[7:3] <= 5)?
                  2
                :
                  2
      :
         (X4[7:2] <= 5)?
           (X6[7:4] <= 7)?
            2
          :
            3
        :
          45
    :
       (X9[7:4] <= 4)?
         (X1[7:4] <= 7)?
          5
        :
          1
      :
         (X5[7:3] <= 7)?
           (X9[7:4] <= 5)?
            13
          :
             (X0[7:4] <= 12)?
               (X9[7:3] <= 9)?
                1
              :
                3
            :
               (X7[7:3] <= 21)?
                1
              :
                2
        :
          2
  :
     (X9[7:4] <= 4)?
       (X10[7:2] <= 31)?
         (X6[7:5] <= 0)?
           (X1[7:3] <= 15)?
             (X3[7:3] <= 3)?
               (X8[7:4] <= 6)?
                 (X7[7:2] <= 30)?
                  5
                :
                   (X8[7:3] <= 11)?
                    1
                  :
                    2
              :
                 (X2[7:3] <= 1)?
                   (X8[7:3] <= 17)?
                    2
                  :
                     (X3[7:2] <= 1)?
                      1
                    :
                      1
                :
                  7
            :
               (X9[7:4] <= 1)?
                 (X1[7:5] <= 3)?
                   (X3[7:1] <= 12)?
                    5
                  :
                     (X0[7:3] <= 8)?
                       (X9[7:4] <= 2)?
                        4
                      :
                        2
                    :
                       (X0[7:5] <= 1)?
                        4
                      :
                         (X8[7:2] <= 28)?
                          6
                        :
                          1
                :
                   (X4[7:4] <= 5)?
                     (X6[7:2] <= 1)?
                      1
                    :
                       (X5[7:4] <= 3)?
                        15
                      :
                        1
                  :
                    1
              :
                 (X4[7:3] <= 5)?
                   (X10[7:3] <= 13)?
                    4
                  :
                     (X0[7:4] <= 6)?
                      1
                    :
                      1
                :
                   (X0[7:5] <= 7)?
                     (X6[7:2] <= 5)?
                      9
                    :
                      1
                  :
                    1
          :
             (X9[7:2] <= 6)?
               (X6[7:4] <= 1)?
                 (X1[7:3] <= 24)?
                   (X1[7:4] <= 7)?
                    1
                  :
                    3
                :
                  2
              :
                1
            :
               (X2[7:4] <= 0)?
                3
              :
                 (X7[7:4] <= 11)?
                  3
                :
                  1
        :
           (X9[7:2] <= 6)?
             (X10[7:2] <= 29)?
               (X3[7:5] <= 2)?
                 (X3[7:3] <= 2)?
                   (X4[7:4] <= 4)?
                    4
                  :
                    8
                :
                  25
              :
                 (X10[7:4] <= 6)?
                  2
                :
                  4
            :
               (X5[7:3] <= 9)?
                 (X2[7:3] <= 3)?
                   (X2[7:3] <= 1)?
                    1
                  :
                    2
                :
                  2
              :
                1
          :
             (X7[7:4] <= 6)?
               (X0[7:3] <= 12)?
                 (X1[7:6] <= 2)?
                   (X10[7:4] <= 4)?
                    1
                  :
                    4
                :
                   (X2[7:1] <= 9)?
                     (X5[7:4] <= 10)?
                       (X0[7:3] <= 11)?
                        19
                      :
                        1
                    :
                      2
                  :
                     (X2[7:4] <= 4)?
                       (X9[7:2] <= 10)?
                        8
                      :
                         (X6[7:3] <= 4)?
                          1
                        :
                          2
                    :
                       (X9[7:2] <= 11)?
                         (X5[7:5] <= 0)?
                           (X3[7:3] <= 5)?
                            4
                          :
                            3
                        :
                          9
                      :
                        2
              :
                 (X0[7:2] <= 23)?
                  1
                :
                  6
            :
              10
      :
         (X1[7:4] <= 5)?
           (X3[7:3] <= 8)?
             (X2[7:1] <= 87)?
               (X0[7:2] <= 0)?
                1
              :
                 (X4[7:2] <= 1)?
                  2
                :
                   (X6[7:5] <= 1)?
                     (X0[7:4] <= 7)?
                       (X0[7:4] <= 5)?
                         (X6[7:2] <= 1)?
                          1
                        :
                           (X6[7:5] <= 1)?
                            9
                          :
                             (X7[7:3] <= 8)?
                              1
                            :
                              1
                      :
                        3
                    :
                      8
                  :
                    20
            :
               (X8[7:3] <= 14)?
                1
              :
                1
          :
             (X2[7:4] <= 8)?
               (X7[7:4] <= 6)?
                1
              :
                2
            :
              5
        :
           (X7[7:2] <= 17)?
             (X8[7:1] <= 107)?
               (X2[7:3] <= 1)?
                 (X9[7:6] <= 1)?
                  3
                :
                  2
              :
                6
            :
              2
          :
             (X1[7:3] <= 14)?
               (X1[7:3] <= 10)?
                1
              :
                 (X4[7:4] <= 1)?
                  1
                :
                  7
            :
               (X1[7:3] <= 14)?
                1
              :
                1
    :
       (X10[7:2] <= 30)?
         (X1[7:3] <= 1)?
           (X6[7:4] <= 5)?
             (X8[7:3] <= 15)?
               (X0[7:3] <= 10)?
                 (X7[7:4] <= 5)?
                   (X10[7:4] <= 8)?
                    1
                  :
                    1
                :
                  2
              :
                 (X2[7:4] <= 10)?
                   (X3[7:4] <= 3)?
                     (X3[7:5] <= 1)?
                       (X6[7:4] <= 0)?
                         (X10[7:3] <= 11)?
                          7
                        :
                           (X1[7:2] <= 7)?
                            1
                          :
                            3
                      :
                         (X0[7:2] <= 26)?
                          3
                        :
                           (X7[7:3] <= 18)?
                             (X7[7:4] <= 7)?
                               (X2[7:2] <= 30)?
                                3
                              :
                                2
                            :
                              11
                          :
                            1
                    :
                       (X8[7:2] <= 19)?
                        1
                      :
                        1
                  :
                    6
                :
                  5
            :
               (X5[7:3] <= 5)?
                 (X9[7:3] <= 9)?
                   (X2[7:3] <= 9)?
                    3
                  :
                     (X2[7:4] <= 9)?
                       (X6[7:2] <= 1)?
                        1
                      :
                         (X6[7:3] <= 1)?
                           (X4[7:4] <= 0)?
                            2
                          :
                            1
                        :
                          2
                    :
                      5
                :
                   (X2[7:3] <= 20)?
                    8
                  :
                    1
              :
                 (X9[7:3] <= 5)?
                  10
                :
                   (X7[7:4] <= 6)?
                    5
                  :
                     (X7[7:3] <= 19)?
                       (X1[7:4] <= 1)?
                         (X10[7:4] <= 2)?
                          2
                        :
                          2
                      :
                        6
                    :
                      2
          :
             (X5[7:3] <= 15)?
               (X2[7:3] <= 18)?
                 (X8[7:3] <= 12)?
                  8
                :
                   (X2[7:3] <= 15)?
                    5
                  :
                    2
              :
                3
            :
               (X0[7:3] <= 10)?
                4
              :
                5
        :
           (X6[7:2] <= 17)?
             (X4[7:4] <= 3)?
               (X1[7:3] <= 13)?
                 (X1[7:1] <= 30)?
                   (X7[7:3] <= 20)?
                     (X7[7:3] <= 17)?
                       (X9[7:4] <= 4)?
                        8
                      :
                         (X7[7:4] <= 3)?
                          2
                        :
                          1
                    :
                      2
                  :
                     (X9[7:2] <= 13)?
                      1
                    :
                      12
                :
                   (X0[7:4] <= 4)?
                     (X8[7:4] <= 12)?
                      17
                    :
                      1
                  :
                     (X1[7:3] <= 7)?
                      3
                    :
                       (X8[7:2] <= 17)?
                        3
                      :
                         (X8[7:4] <= 9)?
                          20
                        :
                           (X2[7:2] <= 5)?
                            6
                          :
                            6
              :
                 (X1[7:4] <= 3)?
                  4
                :
                   (X10[7:5] <= 4)?
                     (X7[7:4] <= 11)?
                      5
                    :
                      3
                  :
                     (X1[7:3] <= 17)?
                      11
                    :
                      1
            :
               (X6[7:2] <= 12)?
                 (X2[7:4] <= 4)?
                   (X3[7:4] <= 1)?
                    2
                  :
                     (X3[7:4] <= 4)?
                       (X3[7:6] <= 1)?
                        4
                      :
                         (X5[7:3] <= 10)?
                          1
                        :
                          1
                    :
                      1
                :
                   (X2[7:4] <= 11)?
                     (X4[7:3] <= 4)?
                      12
                    :
                      1
                  :
                    2
              :
                6
          :
             (X9[7:3] <= 16)?
               (X2[7:3] <= 5)?
                 (X3[7:2] <= 7)?
                  1
                :
                   (X10[7:5] <= 3)?
                    1
                  :
                    1
              :
                15
            :
              4
      :
         (X10[7:4] <= 11)?
           (X9[7:4] <= 3)?
             (X6[7:4] <= 2)?
               (X3[7:4] <= 2)?
                1
              :
                6
            :
               (X3[7:1] <= 9)?
                 (X2[7:3] <= 13)?
                  1
                :
                  1
              :
                 (X0[7:3] <= 21)?
                   (X9[7:4] <= 4)?
                    14
                  :
                    1
                :
                  1
          :
             (X5[7:4] <= 4)?
               (X9[7:3] <= 11)?
                 (X0[7:3] <= 14)?
                  22
                :
                   (X3[7:2] <= 7)?
                    1
                  :
                    3
              :
                 (X5[7:4] <= 2)?
                   (X1[7:2] <= 10)?
                    1
                  :
                    5
                :
                  3
            :
               (X3[7:5] <= 1)?
                 (X10[7:4] <= 10)?
                  4
                :
                   (X2[7:3] <= 0)?
                    3
                  :
                     (X6[7:1] <= 14)?
                      4
                    :
                       (X6[7:4] <= 1)?
                        3
                      :
                         (X4[7:5] <= 0)?
                          2
                        :
                           (X8[7:4] <= 7)?
                             (X10[7:3] <= 19)?
                              2
                            :
                               (X4[7:2] <= 7)?
                                2
                              :
                                1
                          :
                            6
              :
                 (X10[7:4] <= 11)?
                  3
                :
                  1
        :
           (X6[7:2] <= 11)?
             (X4[7:2] <= 6)?
              2
            :
               (X9[7:2] <= 15)?
                3
              :
                2
          :
             (X5[7:4] <= 3)?
              2
            :
              3
;
endmodule
