module top(X0, X1, X2, X3, out);
input [7:0] X0;
input [7:0] X1;
input [7:0] X2;
input [7:0] X3;
output [1:0] out;
assign out = 
   (X0 <= 96)?
     (X2 <= 32)?
       (X1 <= 96)?
         (X3 <= 32)?
          2
        :
           (X0 <= 32)?
            4
          :
             (X3 <= 160)?
               (X1 <= 32)?
                 (X3 <= 96)?
                  1
                :
                  1
              :
                2
            :
               (X3 <= 224)?
                 (X1 <= 32)?
                  1
                :
                  1
              :
                2
      :
         (X3 <= 224)?
           (X3 <= 160)?
            11
          :
             (X0 <= 32)?
               (X1 <= 224)?
                1
              :
                1
            :
              3
        :
           (X1 <= 160)?
            1
          :
            2
    :
       (X3 <= 96)?
         (X1 <= 160)?
           (X2 <= 160)?
             (X0 <= 32)?
               (X3 <= 32)?
                 (X1 <= 32)?
                  1
                :
                  2
              :
                5
            :
               (X1 <= 32)?
                2
              :
                 (X3 <= 32)?
                  3
                :
                   (X2 <= 96)?
                     (X1 <= 96)?
                      1
                    :
                      1
                  :
                     (X1 <= 96)?
                      1
                    :
                      1
          :
             (X3 <= 32)?
               (X0 <= 32)?
                4
              :
                 (X2 <= 224)?
                  1
                :
                  2
            :
              11
        :
           (X2 <= 160)?
             (X0 <= 32)?
               (X3 <= 32)?
                3
              :
                1
            :
              5
          :
             (X3 <= 32)?
               (X0 <= 32)?
                 (X1 <= 224)?
                   (X2 <= 224)?
                    1
                  :
                    1
                :
                   (X2 <= 224)?
                    1
                  :
                    1
              :
                3
            :
               (X0 <= 32)?
                4
              :
                 (X2 <= 224)?
                  1
                :
                   (X1 <= 224)?
                    1
                  :
                    1
      :
         (X1 <= 224)?
          72
        :
           (X2 <= 96)?
             (X0 <= 32)?
              2
            :
               (X3 <= 192)?
                1
              :
                1
          :
            10
  :
     (X3 <= 96)?
       (X1 <= 32)?
         (X2 <= 96)?
           (X0 <= 160)?
             (X2 <= 32)?
              1
            :
              1
          :
            6
        :
           (X3 <= 32)?
             (X0 <= 160)?
              1
            :
               (X2 <= 160)?
                2
              :
                 (X2 <= 224)?
                   (X0 <= 224)?
                    1
                  :
                    1
                :
                  1
          :
            8
      :
         (X2 <= 160)?
          46
        :
           (X3 <= 32)?
            20
          :
             (X1 <= 96)?
               (X0 <= 224)?
                 (X2 <= 224)?
                   (X0 <= 160)?
                    1
                  :
                    1
                :
                  1
              :
                1
            :
               (X0 <= 160)?
                 (X2 <= 224)?
                  3
                :
                  1
              :
                10
    :
       (X2 <= 96)?
         (X1 <= 96)?
           (X2 <= 32)?
             (X1 <= 32)?
               (X0 <= 160)?
                2
              :
                 (X3 <= 160)?
                  2
                :
                   (X0 <= 224)?
                    1
                  :
                     (X3 <= 224)?
                      1
                    :
                      1
            :
              7
          :
             (X1 <= 32)?
              6
            :
               (X3 <= 224)?
                 (X0 <= 160)?
                  1
                :
                   (X0 <= 224)?
                     (X3 <= 160)?
                      1
                    :
                      1
                  :
                    1
              :
                 (X0 <= 224)?
                  2
                :
                  1
        :
           (X0 <= 160)?
             (X3 <= 224)?
              7
            :
               (X2 <= 32)?
                2
              :
                1
          :
            25
      :
         (X1 <= 160)?
           (X0 <= 224)?
             (X1 <= 96)?
              28
            :
               (X3 <= 160)?
                 (X2 <= 224)?
                  2
                :
                  2
              :
                7
          :
             (X2 <= 160)?
               (X3 <= 160)?
                1
              :
                 (X1 <= 96)?
                  2
                :
                  1
            :
              13
        :
           (X2 <= 160)?
             (X0 <= 160)?
               (X3 <= 224)?
                3
              :
                1
            :
              7
          :
             (X3 <= 160)?
               (X0 <= 160)?
                 (X1 <= 224)?
                   (X2 <= 224)?
                    1
                  :
                    1
                :
                  1
              :
                6
            :
               (X0 <= 160)?
                6
              :
                 (X2 <= 224)?
                   (X1 <= 224)?
                     (X3 <= 224)?
                       (X0 <= 224)?
                        1
                      :
                        1
                    :
                       (X0 <= 224)?
                        1
                      :
                        1
                  :
                    2
                :
                   (X3 <= 224)?
                     (X0 <= 224)?
                      1
                    :
                      1
                  :
                    2
;
endmodule
