module top(X13, X27, X235, X264, X278, out);
input [7:0] X13;
input [7:0] X27;
input [7:0] X235;
input [7:0] X264;
input [7:0] X278;
output [4:0] out;
assign out = 
   (X278[7:6] <= 0)?
    167
  :
     (X278[7:5] <= 1)?
      24
    :
       (X278[7:3] <= 15)?
         (X13[7:5] <= 1)?
           (X27[7:6] <= 4)?
            17
          :
            1
        :
           (X278[7:4] <= 3)?
            11
          :
             (X278[7:6] <= 1)?
              7
            :
               (X278[7:5] <= 7)?
                9
              :
                 (X235[7:6] <= 4)?
                   (X264[7:4] <= 7)?
                    2
                  :
                    1
                :
                  6
      :
         (X278[7:4] <= 15)?
          33
        :
           (X278[7:6] <= 1)?
            4
          :
            12
;
endmodule
