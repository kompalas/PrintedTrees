module top(X0, X1, X2, X3, X4, X5, X6, X7, X8, X9, X10, out);
input [7:0] X0;
input [7:0] X1;
input [7:0] X2;
input [7:0] X3;
input [7:0] X4;
input [7:0] X5;
input [7:0] X6;
input [7:0] X7;
input [7:0] X8;
input [7:0] X9;
input [7:0] X10;
output [3:0] out;
assign out = 
   (X10 <= 84)?
     (X9 <= 31)?
       (X1 <= 132)?
         (X1 <= 66)?
           (X4 <= 30)?
             (X1 <= 40)?
               (X4 <= 18)?
                1
              :
                6
            :
               (X6 <= 26)?
                 (X5 <= 27)?
                   (X4 <= 27)?
                    2
                  :
                    1
                :
                  3
              :
                 (X0 <= 46)?
                  1
                :
                  7
          :
             (X10 <= 69)?
              19
            :
               (X5 <= 36)?
                2
              :
                2
        :
           (X6 <= 56)?
             (X10 <= 77)?
               (X2 <= 29)?
                 (X6 <= 6)?
                   (X7 <= 120)?
                    5
                  :
                    1
                :
                  33
              :
                 (X2 <= 49)?
                  2
                :
                   (X4 <= 18)?
                    2
                  :
                     (X8 <= 99)?
                      11
                    :
                       (X4 <= 29)?
                        4
                      :
                         (X8 <= 123)?
                           (X6 <= 53)?
                            4
                          :
                            1
                        :
                          2
            :
               (X6 <= 12)?
                1
              :
                1
          :
             (X7 <= 121)?
               (X8 <= 80)?
                1
              :
                22
            :
               (X4 <= 36)?
                 (X3 <= 26)?
                  3
                :
                   (X3 <= 49)?
                    5
                  :
                     (X9 <= 25)?
                      1
                    :
                      4
              :
                6
      :
         (X3 <= 17)?
          4
        :
           (X1 <= 133)?
            1
          :
             (X1 <= 144)?
               (X6 <= 71)?
                1
              :
                1
            :
              7
    :
       (X6 <= 68)?
         (X1 <= 80)?
           (X9 <= 51)?
             (X2 <= 81)?
               (X0 <= 89)?
                 (X2 <= 22)?
                   (X6 <= 37)?
                     (X4 <= 26)?
                       (X10 <= 59)?
                        5
                      :
                         (X0 <= 80)?
                          2
                        :
                          1
                    :
                      10
                  :
                    1
                :
                   (X4 <= 24)?
                     (X7 <= 107)?
                      1
                    :
                      5
                  :
                     (X2 <= 42)?
                       (X3 <= 22)?
                         (X4 <= 30)?
                          8
                        :
                          1
                      :
                         (X7 <= 129)?
                           (X7 <= 111)?
                            3
                          :
                             (X1 <= 55)?
                              2
                            :
                              2
                        :
                          4
                    :
                       (X10 <= 28)?
                        4
                      :
                         (X1 <= 38)?
                          2
                        :
                           (X3 <= 15)?
                            4
                          :
                             (X4 <= 31)?
                               (X4 <= 29)?
                                 (X3 <= 18)?
                                  5
                                :
                                   (X9 <= 36)?
                                     (X1 <= 57)?
                                      4
                                    :
                                       (X3 <= 28)?
                                        2
                                      :
                                        1
                                  :
                                     (X8 <= 116)?
                                      1
                                    :
                                      6
                              :
                                4
                            :
                              4
              :
                11
            :
               (X5 <= 25)?
                 (X1 <= 62)?
                   (X1 <= 52)?
                     (X3 <= 22)?
                      4
                    :
                       (X1 <= 48)?
                        4
                      :
                        1
                  :
                    5
                :
                  5
              :
                 (X9 <= 41)?
                   (X3 <= 24)?
                     (X7 <= 139)?
                       (X7 <= 124)?
                         (X9 <= 34)?
                          1
                        :
                          2
                      :
                        5
                    :
                      3
                  :
                    6
                :
                   (X7 <= 143)?
                     (X8 <= 114)?
                      2
                    :
                      1
                  :
                     (X1 <= 53)?
                      9
                    :
                       (X6 <= 28)?
                        1
                      :
                        2
          :
             (X4 <= 49)?
               (X10 <= 49)?
                 (X7 <= 124)?
                  6
                :
                   (X6 <= 9)?
                     (X2 <= 170)?
                      4
                    :
                      1
                  :
                     (X0 <= 216)?
                      22
                    :
                      1
              :
                 (X8 <= 57)?
                   (X6 <= 26)?
                     (X0 <= 180)?
                      1
                    :
                      1
                  :
                    2
                :
                   (X9 <= 105)?
                     (X1 <= 50)?
                       (X10 <= 81)?
                         (X2 <= 109)?
                           (X10 <= 61)?
                             (X3 <= 20)?
                              3
                            :
                               (X1 <= 44)?
                                1
                              :
                                1
                          :
                             (X1 <= 22)?
                              3
                            :
                               (X3 <= 29)?
                                3
                              :
                                2
                        :
                           (X6 <= 5)?
                            1
                          :
                             (X3 <= 47)?
                              16
                            :
                              1
                      :
                         (X3 <= 29)?
                          1
                        :
                          3
                    :
                       (X4 <= 38)?
                        16
                      :
                        1
                  :
                     (X3 <= 19)?
                      1
                    :
                      1
            :
               (X7 <= 151)?
                 (X6 <= 5)?
                  1
                :
                   (X9 <= 122)?
                     (X9 <= 82)?
                      3
                    :
                      4
                  :
                    4
              :
                 (X1 <= 59)?
                  1
                :
                  2
        :
           (X10 <= 62)?
             (X10 <= 26)?
               (X8 <= 110)?
                2
              :
                5
            :
               (X1 <= 111)?
                 (X7 <= 118)?
                  10
                :
                   (X0 <= 48)?
                    7
                  :
                     (X6 <= 61)?
                       (X8 <= 114)?
                         (X7 <= 185)?
                           (X4 <= 26)?
                             (X4 <= 24)?
                              2
                            :
                              2
                          :
                             (X2 <= 35)?
                               (X4 <= 34)?
                                7
                              :
                                2
                            :
                              13
                        :
                          3
                      :
                         (X6 <= 18)?
                           (X0 <= 92)?
                            11
                          :
                            1
                        :
                           (X1 <= 99)?
                             (X2 <= 1)?
                              4
                            :
                               (X2 <= 17)?
                                8
                              :
                                 (X2 <= 44)?
                                   (X4 <= 37)?
                                    6
                                  :
                                    1
                                :
                                  3
                          :
                            9
                    :
                       (X6 <= 63)?
                        1
                      :
                        4
              :
                 (X7 <= 157)?
                   (X1 <= 144)?
                     (X6 <= 10)?
                       (X8 <= 121)?
                        1
                      :
                         (X6 <= 5)?
                          1
                        :
                          1
                    :
                      9
                  :
                     (X5 <= 41)?
                      1
                    :
                       (X8 <= 106)?
                        1
                      :
                        1
                :
                   (X10 <= 47)?
                    3
                  :
                    1
          :
             (X9 <= 48)?
               (X3 <= 11)?
                2
              :
                 (X9 <= 33)?
                  5
                :
                   (X1 <= 85)?
                     (X9 <= 44)?
                       (X6 <= 13)?
                         (X2 <= 70)?
                          1
                        :
                          1
                      :
                        6
                    :
                       (X8 <= 155)?
                        5
                      :
                        1
                  :
                     (X5 <= 31)?
                       (X1 <= 96)?
                        4
                      :
                         (X9 <= 38)?
                          1
                        :
                          4
                    :
                      13
            :
               (X5 <= 23)?
                 (X6 <= 36)?
                   (X4 <= 29)?
                     (X9 <= 74)?
                      1
                    :
                      1
                  :
                    4
                :
                  2
              :
                 (X6 <= 13)?
                  1
                :
                  9
      :
         (X6 <= 91)?
           (X2 <= 116)?
             (X5 <= 153)?
               (X5 <= 92)?
                 (X9 <= 103)?
                   (X5 <= 49)?
                    10
                  :
                     (X1 <= 63)?
                      3
                    :
                       (X7 <= 115)?
                         (X8 <= 122)?
                          4
                        :
                          1
                      :
                         (X1 <= 92)?
                           (X3 <= 29)?
                             (X9 <= 36)?
                              2
                            :
                              3
                          :
                            4
                        :
                          6
                :
                  2
              :
                8
            :
              2
          :
             (X0 <= 69)?
              1
            :
              6
        :
           (X10 <= 30)?
            1
          :
             (X8 <= 98)?
               (X4 <= 26)?
                1
              :
                 (X10 <= 57)?
                  13
                :
                  1
            :
              26
  :
     (X1 <= 57)?
       (X10 <= 124)?
         (X8 <= 104)?
           (X1 <= 45)?
             (X1 <= 39)?
               (X0 <= 133)?
                 (X7 <= 96)?
                   (X7 <= 73)?
                    1
                  :
                    4
                :
                   (X8 <= 98)?
                    7
                  :
                    3
              :
                8
            :
               (X9 <= 58)?
                2
              :
                5
          :
             (X8 <= 79)?
              8
            :
               (X8 <= 93)?
                 (X3 <= 16)?
                  1
                :
                   (X4 <= 38)?
                     (X8 <= 87)?
                       (X3 <= 20)?
                        1
                      :
                        2
                    :
                      1
                  :
                    1
              :
                5
        :
           (X10 <= 116)?
             (X0 <= 157)?
               (X4 <= 27)?
                 (X2 <= 120)?
                   (X3 <= 15)?
                    3
                  :
                     (X2 <= 42)?
                      2
                    :
                       (X1 <= 14)?
                        2
                      :
                         (X2 <= 69)?
                          2
                        :
                          7
                :
                   (X5 <= 16)?
                    1
                  :
                    7
              :
                 (X7 <= 150)?
                   (X6 <= 78)?
                     (X9 <= 55)?
                       (X4 <= 32)?
                         (X0 <= 62)?
                          1
                        :
                          3
                      :
                        4
                    :
                      8
                  :
                    2
                :
                   (X10 <= 106)?
                    4
                  :
                    1
            :
              2
          :
             (X0 <= 56)?
               (X2 <= 31)?
                1
              :
                2
            :
              7
      :
         (X3 <= 66)?
           (X9 <= 61)?
             (X6 <= 8)?
               (X7 <= 86)?
                8
              :
                 (X7 <= 110)?
                   (X8 <= 115)?
                    4
                  :
                    1
                :
                  3
            :
               (X3 <= 18)?
                 (X0 <= 100)?
                  9
                :
                  2
              :
                 (X5 <= 72)?
                   (X3 <= 28)?
                    13
                  :
                     (X3 <= 31)?
                      2
                    :
                       (X10 <= 146)?
                         (X8 <= 98)?
                          2
                        :
                          2
                      :
                        4
                :
                   (X0 <= 14)?
                    1
                  :
                    4
          :
             (X6 <= 37)?
               (X8 <= 100)?
                 (X5 <= 23)?
                  2
                :
                  3
              :
                 (X0 <= 71)?
                   (X9 <= 74)?
                    4
                  :
                     (X6 <= 28)?
                      3
                    :
                      1
                :
                  20
            :
               (X0 <= 12)?
                 (X8 <= 194)?
                  1
                :
                  1
              :
                5
        :
           (X8 <= 51)?
            1
          :
             (X5 <= 11)?
               (X10 <= 134)?
                1
              :
                1
            :
              8
    :
       (X9 <= 39)?
         (X1 <= 154)?
           (X5 <= 92)?
             (X2 <= 24)?
               (X3 <= 24)?
                 (X1 <= 73)?
                   (X5 <= 54)?
                    1
                  :
                    1
                :
                   (X9 <= 38)?
                    11
                  :
                    1
              :
                 (X10 <= 96)?
                   (X7 <= 120)?
                     (X2 <= 1)?
                      4
                    :
                      2
                  :
                    4
                :
                   (X3 <= 51)?
                    5
                  :
                     (X9 <= 19)?
                      1
                    :
                      2
            :
               (X2 <= 82)?
                11
              :
                 (X4 <= 30)?
                  2
                :
                  3
          :
             (X8 <= 147)?
              6
            :
               (X8 <= 158)?
                2
              :
                 (X6 <= 42)?
                  1
                :
                  1
        :
           (X4 <= 31)?
             (X5 <= 32)?
              1
            :
              2
          :
            3
      :
         (X10 <= 175)?
           (X4 <= 35)?
             (X3 <= 71)?
               (X4 <= 24)?
                 (X2 <= 12)?
                   (X10 <= 124)?
                    5
                  :
                     (X0 <= 12)?
                      2
                    :
                      4
                :
                   (X3 <= 27)?
                     (X1 <= 76)?
                       (X3 <= 24)?
                        5
                      :
                        1
                    :
                       (X4 <= 16)?
                         (X0 <= 37)?
                          2
                        :
                          1
                      :
                        5
                  :
                     (X9 <= 51)?
                      4
                    :
                      2
              :
                 (X3 <= 25)?
                   (X10 <= 167)?
                    35
                  :
                    1
                :
                   (X9 <= 54)?
                     (X1 <= 86)?
                      13
                    :
                       (X6 <= 16)?
                        4
                      :
                         (X2 <= 1)?
                          1
                        :
                          3
                  :
                     (X8 <= 108)?
                      5
                    :
                       (X8 <= 136)?
                         (X5 <= 41)?
                          1
                        :
                          6
                      :
                         (X8 <= 167)?
                          5
                        :
                          2
            :
              3
          :
             (X10 <= 112)?
               (X4 <= 45)?
                7
              :
                 (X10 <= 100)?
                  4
                :
                   (X5 <= 34)?
                    2
                  :
                    1
            :
               (X2 <= 131)?
                 (X5 <= 40)?
                   (X8 <= 121)?
                    1
                  :
                    2
                :
                  5
              :
                 (X9 <= 90)?
                  4
                :
                  2
        :
           (X6 <= 75)?
             (X7 <= 61)?
              3
            :
               (X9 <= 63)?
                1
              :
                3
          :
             (X9 <= 64)?
              1
            :
              2
;
endmodule
