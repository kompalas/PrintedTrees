module dt(X13, X186, X219, X278, out);
input [7:0] X13;
input [7:0] X186;
input [7:0] X219;
input [7:0] X278;
output [4:0] out;
assign out = 
   (X278 <= 8)?
    172
  :
     (X278 <= 24)?
      22
    :
       (X278 <= 136)?
         (X13 <= 24)?
           (X219 <= 64)?
            1
          :
            19
        :
           (X278 <= 40)?
            8
          :
             (X278 <= 56)?
              9
            :
               (X13 <= 80)?
                 (X278 <= 120)?
                   (X186 <= 80)?
                    1
                  :
                    1
                :
                  7
              :
                7
      :
         (X278 <= 176)?
          31
        :
           (X278 <= 232)?
            2
          :
            14
;
endmodule
