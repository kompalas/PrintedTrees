module top(X0, X1, X2, X3, X4, X5, X6, X7, X8, X9, X10, out);
input [7:0] X0;
input [7:0] X1;
input [7:0] X2;
input [7:0] X3;
input [7:0] X4;
input [7:0] X5;
input [7:0] X6;
input [7:0] X7;
input [7:0] X8;
input [7:0] X9;
input [7:0] X10;
output [3:0] out;
assign out = 
   (X10[7:3] <= 11)?
     (X0[7:1] <= 70)?
       (X6[7:3] <= 11)?
         (X9[7:2] <= 6)?
           (X3[7:4] <= 7)?
             (X4[7:4] <= 2)?
               (X6[7:1] <= 40)?
                 (X2[7:3] <= 11)?
                   (X9[7:3] <= 4)?
                     (X0[7:4] <= 6)?
                       (X9[7:5] <= 3)?
                        13
                      :
                         (X0[7:4] <= 4)?
                           (X4[7:2] <= 7)?
                            1
                          :
                            5
                        :
                          2
                    :
                       (X10[7:4] <= 5)?
                        1
                      :
                        2
                  :
                    20
                :
                   (X1[7:3] <= 3)?
                    1
                  :
                     (X9[7:2] <= 9)?
                      1
                    :
                      4
              :
                3
            :
               (X4[7:3] <= 9)?
                 (X7[7:3] <= 18)?
                  20
                :
                   (X7[7:2] <= 36)?
                     (X0[7:2] <= 19)?
                      2
                    :
                      3
                  :
                    12
              :
                1
          :
             (X2[7:3] <= 7)?
              1
            :
              3
        :
           (X1[7:1] <= 47)?
             (X1[7:3] <= 3)?
              5
            :
               (X0[7:3] <= 12)?
                 (X1[7:1] <= 23)?
                   (X7[7:2] <= 29)?
                    3
                  :
                     (X6[7:4] <= 7)?
                       (X1[7:2] <= 11)?
                        7
                      :
                         (X10[7:3] <= 11)?
                          1
                        :
                          1
                    :
                      1
                :
                   (X0[7:1] <= 24)?
                    11
                  :
                     (X2[7:2] <= 0)?
                      8
                    :
                       (X6[7:1] <= 17)?
                         (X7[7:3] <= 15)?
                          7
                        :
                           (X7[7:1] <= 72)?
                             (X0[7:1] <= 41)?
                               (X4[7:3] <= 11)?
                                 (X8[7:2] <= 31)?
                                  11
                                :
                                   (X8[7:4] <= 10)?
                                    3
                                  :
                                     (X10[7:3] <= 8)?
                                      1
                                    :
                                       (X9[7:2] <= 13)?
                                        1
                                      :
                                        7
                              :
                                2
                            :
                              3
                          :
                             (X8[7:3] <= 15)?
                               (X7[7:3] <= 21)?
                                1
                              :
                                1
                            :
                              8
                      :
                         (X3[7:5] <= 3)?
                          14
                        :
                           (X0[7:3] <= 10)?
                             (X4[7:2] <= 9)?
                               (X4[7:3] <= 2)?
                                 (X1[7:2] <= 13)?
                                  1
                                :
                                  13
                              :
                                 (X1[7:3] <= 10)?
                                   (X2[7:4] <= 7)?
                                     (X1[7:3] <= 7)?
                                      2
                                    :
                                       (X0[7:4] <= 6)?
                                        3
                                      :
                                        1
                                  :
                                    4
                                :
                                  7
                            :
                              10
                          :
                             (X9[7:3] <= 6)?
                              1
                            :
                              8
              :
                 (X0[7:2] <= 31)?
                   (X9[7:2] <= 15)?
                     (X9[7:2] <= 12)?
                      18
                    :
                       (X0[7:3] <= 17)?
                        1
                      :
                        1
                  :
                     (X0[7:3] <= 13)?
                       (X9[7:2] <= 13)?
                        3
                      :
                         (X9[7:2] <= 41)?
                          7
                        :
                          1
                    :
                       (X7[7:1] <= 103)?
                        13
                      :
                         (X1[7:1] <= 37)?
                          1
                        :
                          2
                :
                   (X2[7:1] <= 65)?
                     (X0[7:1] <= 70)?
                      7
                    :
                      1
                  :
                    5
          :
             (X10[7:3] <= 3)?
              2
            :
               (X1[7:3] <= 16)?
                 (X0[7:3] <= 11)?
                   (X8[7:2] <= 23)?
                     (X5[7:2] <= 9)?
                       (X10[7:5] <= 2)?
                        2
                      :
                        1
                    :
                      8
                  :
                     (X7[7:5] <= 4)?
                       (X9[7:2] <= 7)?
                         (X5[7:2] <= 8)?
                          2
                        :
                          3
                      :
                         (X0[7:2] <= 15)?
                           (X4[7:4] <= 6)?
                             (X7[7:5] <= 5)?
                              6
                            :
                              1
                          :
                            2
                        :
                          13
                    :
                      13
                :
                   (X10[7:4] <= 3)?
                    3
                  :
                     (X2[7:2] <= 7)?
                      1
                    :
                      1
              :
                 (X9[7:3] <= 9)?
                  2
                :
                  2
      :
         (X4[7:3] <= 2)?
           (X6[7:3] <= 17)?
            2
          :
            3
        :
          45
    :
       (X9[7:3] <= 6)?
         (X1[7:4] <= 5)?
          5
        :
          1
      :
         (X5[7:1] <= 34)?
           (X9[7:3] <= 9)?
            13
          :
             (X0[7:3] <= 24)?
               (X9[7:2] <= 18)?
                1
              :
                3
            :
               (X7[7:4] <= 13)?
                1
              :
                2
        :
          2
  :
     (X9[7:3] <= 7)?
       (X10[7:2] <= 32)?
         (X6[7:5] <= 0)?
           (X1[7:1] <= 56)?
             (X3[7:3] <= 4)?
               (X8[7:5] <= 3)?
                 (X7[7:3] <= 17)?
                  5
                :
                   (X8[7:2] <= 19)?
                    1
                  :
                    2
              :
                 (X2[7:3] <= 1)?
                   (X8[7:3] <= 18)?
                    2
                  :
                     (X3[7:1] <= 6)?
                      1
                    :
                      1
                :
                  7
            :
               (X9[7:2] <= 10)?
                 (X1[7:4] <= 5)?
                   (X3[7:2] <= 6)?
                    5
                  :
                     (X0[7:3] <= 8)?
                       (X9[7:2] <= 12)?
                        4
                      :
                        2
                    :
                       (X0[7:4] <= 4)?
                        4
                      :
                         (X8[7:4] <= 10)?
                          6
                        :
                          1
                :
                   (X4[7:5] <= 3)?
                     (X6[7:3] <= 0)?
                      1
                    :
                       (X5[7:1] <= 24)?
                        15
                      :
                        1
                  :
                    1
              :
                 (X4[7:3] <= 5)?
                   (X10[7:2] <= 24)?
                    4
                  :
                     (X0[7:4] <= 6)?
                      1
                    :
                      1
                :
                   (X0[7:3] <= 17)?
                     (X6[7:1] <= 11)?
                      9
                    :
                      1
                  :
                    1
          :
             (X9[7:3] <= 4)?
               (X6[7:4] <= 1)?
                 (X1[7:3] <= 21)?
                   (X1[7:2] <= 33)?
                    1
                  :
                    3
                :
                  2
              :
                1
            :
               (X2 <= 6)?
                3
              :
                 (X7[7:3] <= 18)?
                  3
                :
                  1
        :
           (X9[7:2] <= 9)?
             (X10[7:3] <= 16)?
               (X3[7:3] <= 6)?
                 (X3[7:2] <= 7)?
                   (X4[7:3] <= 5)?
                    4
                  :
                    8
                :
                  25
              :
                 (X10[7:1] <= 34)?
                  2
                :
                  4
            :
               (X5[7:2] <= 21)?
                 (X2[7:3] <= 3)?
                   (X2[7:3] <= 1)?
                    1
                  :
                    2
                :
                  2
              :
                1
          :
             (X7[7:2] <= 39)?
               (X0[7:3] <= 13)?
                 (X1[7:4] <= 3)?
                   (X10[7:1] <= 33)?
                    1
                  :
                    4
                :
                   (X2[7:1] <= 9)?
                     (X5[7:2] <= 32)?
                       (X0[7:3] <= 9)?
                        19
                      :
                        1
                    :
                      2
                  :
                     (X2[7:3] <= 8)?
                       (X9[7:1] <= 20)?
                        8
                      :
                         (X6[7:3] <= 5)?
                          1
                        :
                          2
                    :
                       (X9 <= 44)?
                         (X5[7:1] <= 28)?
                           (X3[7:3] <= 6)?
                            4
                          :
                            3
                        :
                          9
                      :
                        2
              :
                 (X0[7:2] <= 23)?
                  1
                :
                  6
            :
              10
      :
         (X1[7:3] <= 10)?
           (X3[7:3] <= 11)?
             (X2[7:1] <= 88)?
               (X0[7:2] <= 4)?
                1
              :
                 (X4[7:3] <= 2)?
                  2
                :
                   (X6[7:4] <= 1)?
                     (X0[7:3] <= 15)?
                       (X0[7:3] <= 11)?
                         (X6[7:2] <= 2)?
                          1
                        :
                           (X6[7:5] <= 2)?
                            9
                          :
                             (X7[7:4] <= 8)?
                              1
                            :
                              1
                      :
                        3
                    :
                      8
                  :
                    20
            :
               (X8[7:3] <= 13)?
                1
              :
                1
          :
             (X2[7:4] <= 7)?
               (X7[7:3] <= 17)?
                1
              :
                2
            :
              5
        :
           (X7[7:3] <= 9)?
             (X8[7:3] <= 27)?
               (X2[7:3] <= 1)?
                 (X9[7:3] <= 5)?
                  3
                :
                  2
              :
                6
            :
              2
          :
             (X1[7:3] <= 15)?
               (X1[7:3] <= 10)?
                1
              :
                 (X4[7:3] <= 4)?
                  1
                :
                  7
            :
               (X1[7:3] <= 15)?
                1
              :
                1
    :
       (X10[7:2] <= 31)?
         (X1[7:3] <= 5)?
           (X6[7:3] <= 8)?
             (X8[7:3] <= 15)?
               (X0[7:3] <= 9)?
                 (X7[7:4] <= 5)?
                   (X10[7:3] <= 18)?
                    1
                  :
                    1
                :
                  2
              :
                 (X2[7:2] <= 42)?
                   (X3[7:3] <= 5)?
                     (X3[7:4] <= 3)?
                       (X6[7:4] <= 1)?
                         (X10[7:2] <= 21)?
                          7
                        :
                           (X1[7:2] <= 7)?
                            1
                          :
                            3
                      :
                         (X0[7:3] <= 12)?
                          3
                        :
                           (X7[7:1] <= 83)?
                             (X7[7:4] <= 7)?
                               (X2[7:2] <= 30)?
                                3
                              :
                                2
                            :
                              11
                          :
                            1
                    :
                       (X8[7:2] <= 19)?
                        1
                      :
                        1
                  :
                    6
                :
                  5
            :
               (X5[7:2] <= 9)?
                 (X9[7:3] <= 9)?
                   (X2[7:2] <= 28)?
                    3
                  :
                     (X2[7:2] <= 30)?
                       (X6[7:2] <= 1)?
                        1
                      :
                         (X6[7:1] <= 8)?
                           (X4[7:2] <= 8)?
                            2
                          :
                            1
                        :
                          2
                    :
                      5
                :
                   (X2[7:3] <= 20)?
                    8
                  :
                    1
              :
                 (X9[7:4] <= 8)?
                  10
                :
                   (X7[7:3] <= 17)?
                    5
                  :
                     (X7[7:2] <= 38)?
                       (X1[7:3] <= 5)?
                         (X10[7:2] <= 23)?
                          2
                        :
                          2
                      :
                        6
                    :
                      2
          :
             (X5[7:2] <= 33)?
               (X2[7:3] <= 18)?
                 (X8[7:2] <= 31)?
                  8
                :
                   (X2[7:2] <= 29)?
                    5
                  :
                    2
              :
                3
            :
               (X0[7:2] <= 25)?
                4
              :
                5
        :
           (X6[7:2] <= 18)?
             (X4[7:2] <= 12)?
               (X1[7:2] <= 23)?
                 (X1[7:1] <= 32)?
                   (X7[7:1] <= 67)?
                     (X7[7:3] <= 17)?
                       (X9[7:4] <= 7)?
                        8
                      :
                         (X7[7:2] <= 24)?
                          2
                        :
                          1
                    :
                      2
                  :
                     (X9[7:3] <= 7)?
                      1
                    :
                      12
                :
                   (X0[7:5] <= 5)?
                     (X8[7:4] <= 12)?
                      17
                    :
                      1
                  :
                     (X1[7:3] <= 7)?
                      3
                    :
                       (X8[7:4] <= 7)?
                        3
                      :
                         (X8[7:3] <= 15)?
                          20
                        :
                           (X2[7:3] <= 2)?
                            6
                          :
                            6
              :
                 (X1[7:5] <= 3)?
                  4
                :
                   (X10[7:4] <= 7)?
                     (X7[7:3] <= 21)?
                      5
                    :
                      3
                  :
                     (X1[7:1] <= 69)?
                      11
                    :
                      1
            :
               (X6[7:1] <= 25)?
                 (X2[7:4] <= 4)?
                   (X3[7:4] <= 2)?
                    2
                  :
                     (X3[7:2] <= 14)?
                       (X3 <= 35)?
                        4
                      :
                         (X5[7:3] <= 10)?
                          1
                        :
                          1
                    :
                      1
                :
                   (X2[7:2] <= 39)?
                     (X4[7:4] <= 4)?
                      12
                    :
                      1
                  :
                    2
              :
                6
          :
             (X9[7:2] <= 35)?
               (X2[7:3] <= 8)?
                 (X3[7:3] <= 6)?
                  1
                :
                   (X10[7:4] <= 9)?
                    1
                  :
                    1
              :
                15
            :
              4
      :
         (X10[7:2] <= 46)?
           (X9 <= 56)?
             (X6[7:4] <= 3)?
               (X3[7:4] <= 1)?
                1
              :
                6
            :
               (X3[7:1] <= 11)?
                 (X2[7:1] <= 55)?
                  1
                :
                  1
              :
                 (X0[7:4] <= 16)?
                   (X9[7:4] <= 4)?
                    14
                  :
                    1
                :
                  1
          :
             (X5[7:2] <= 14)?
               (X9[7:3] <= 11)?
                 (X0[7:4] <= 7)?
                  22
                :
                   (X3[7:2] <= 8)?
                    1
                  :
                    3
              :
                 (X5[7:4] <= 2)?
                   (X1[7:5] <= 2)?
                    1
                  :
                    5
                :
                  3
            :
               (X3[7:5] <= 1)?
                 (X10[7:5] <= 6)?
                  4
                :
                   (X2[7:1] <= 6)?
                    3
                  :
                     (X6[7:1] <= 13)?
                      4
                    :
                       (X6[7:2] <= 9)?
                        3
                      :
                         (X4[7:4] <= 1)?
                          2
                        :
                           (X8[7:4] <= 8)?
                             (X10[7:4] <= 11)?
                              2
                            :
                               (X4[7:1] <= 12)?
                                2
                              :
                                1
                          :
                            6
              :
                 (X10[7:4] <= 11)?
                  3
                :
                  1
        :
           (X6[7:3] <= 7)?
             (X4[7:2] <= 7)?
              2
            :
               (X9[7:2] <= 17)?
                3
              :
                2
          :
             (X5[7:1] <= 41)?
              2
            :
              3
;
endmodule
