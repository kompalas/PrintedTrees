module top(X0, X1, X2, X3, X4, out);
input [7:0] X0;
input [7:0] X1;
input [7:0] X2;
input [7:0] X3;
input [7:0] X4;
output [0:0] out;
assign out = 
   (X0[7:6] <= 0)?
     (X2[7:6] <= 0)?
       (X1[7:6] <= 0)?
         (X3[7:6] <= 1)?
           (X4[7:6] <= 0)?
            1
          :
             (X1[7:5] <= 0)?
              42
            :
               (X1[7:6] <= 0)?
                 (X4[7:6] <= 0)?
                  17
                :
                   (X1[7:6] <= 0)?
                     (X1[7:6] <= 0)?
                       (X1[7:6] <= 0)?
                         (X1[7:6] <= 0)?
                           (X2[7:6] <= 0)?
                            3
                          :
                            2
                        :
                          17
                      :
                         (X0[7:6] <= 0)?
                          3
                        :
                           (X3[7:6] <= 0)?
                             (X1[7:6] <= 0)?
                               (X2[7:6] <= 0)?
                                3
                              :
                                4
                            :
                               (X2[7:6] <= 0)?
                                 (X1[7:6] <= 1)?
                                  2
                                :
                                  3
                              :
                                2
                          :
                            2
                    :
                       (X1[7:5] <= 1)?
                        40
                      :
                         (X1[7:6] <= 0)?
                           (X2[7:6] <= 0)?
                             (X1[7:6] <= 0)?
                              1
                            :
                              6
                          :
                            4
                        :
                          12
                  :
                     (X2[7:6] <= 0)?
                      2
                    :
                      1
              :
                22
        :
           (X1[7:6] <= 0)?
            5
          :
             (X3[7:6] <= 2)?
               (X2[7:5] <= 0)?
                1
              :
                 (X1[7:5] <= 0)?
                   (X1[7:5] <= 1)?
                    1
                  :
                    2
                :
                   (X1[7:6] <= 0)?
                     (X1[7:5] <= 1)?
                      1
                    :
                      1
                  :
                    2
            :
              1
      :
         (X1[7:6] <= 0)?
           (X1[7:6] <= 1)?
             (X2[7:6] <= 0)?
               (X4[7:6] <= 0)?
                1
              :
                 (X3[7:6] <= 0)?
                   (X3[7:4] <= 0)?
                     (X1[7:5] <= 3)?
                       (X1[7:6] <= 0)?
                        1
                      :
                         (X0[7:5] <= 0)?
                          1
                        :
                           (X1[7:6] <= 0)?
                            1
                          :
                            2
                    :
                      1
                  :
                    1
                :
                  1
            :
               (X3[7:6] <= 0)?
                5
              :
                1
          :
            2
        :
           (X4[7:5] <= 0)?
             (X1[7:5] <= 3)?
              1
            :
              1
          :
            9
    :
       (X1[7:5] <= 3)?
         (X1[7:6] <= 0)?
           (X1[7:6] <= 0)?
             (X1[7:6] <= 0)?
              2
            :
               (X1[7:6] <= 0)?
                1
              :
                 (X1[7:5] <= 3)?
                   (X1[7:6] <= 0)?
                     (X1[7:6] <= 1)?
                       (X3[7:5] <= 3)?
                        6
                      :
                        1
                    :
                       (X0[7:6] <= 0)?
                        1
                      :
                         (X3[7:6] <= 0)?
                           (X1[7:6] <= 0)?
                             (X3[7:4] <= 7)?
                               (X3[7:6] <= 0)?
                                 (X1[7:5] <= 2)?
                                  2
                                :
                                  2
                              :
                                 (X1[7:4] <= 2)?
                                  2
                                :
                                  1
                            :
                               (X1[7:6] <= 0)?
                                 (X4[7:6] <= 0)?
                                  1
                                :
                                  1
                              :
                                3
                          :
                            2
                        :
                          1
                  :
                     (X3[7:5] <= 3)?
                      6
                    :
                      1
                :
                   (X2[7:6] <= 1)?
                    1
                  :
                    2
          :
            6
        :
           (X1[7:6] <= 0)?
             (X1[7:5] <= 0)?
               (X4[7:5] <= 3)?
                 (X1[7:6] <= 1)?
                  1
                :
                   (X2[7:6] <= 0)?
                    1
                  :
                     (X3[7:6] <= 0)?
                      1
                    :
                      1
              :
                1
            :
               (X1[7:4] <= 5)?
                 (X3[7:5] <= 4)?
                  3
                :
                   (X1[7:5] <= 4)?
                    1
                  :
                     (X3[7:6] <= 3)?
                       (X2[7:4] <= 10)?
                        1
                      :
                        1
                    :
                      2
              :
                 (X3[7:6] <= 0)?
                  1
                :
                   (X4[7:6] <= 1)?
                    1
                  :
                     (X0[7:6] <= 0)?
                      1
                    :
                       (X3[7:6] <= 0)?
                         (X1[7:5] <= 1)?
                           (X3[7:6] <= 0)?
                            2
                          :
                             (X1[7:5] <= 1)?
                               (X2[7:6] <= 1)?
                                1
                              :
                                1
                            :
                              2
                        :
                           (X2[7:5] <= 5)?
                            2
                          :
                             (X1[7:6] <= 0)?
                               (X3[7:5] <= 1)?
                                1
                              :
                                1
                            :
                              1
                      :
                         (X1[7:5] <= 1)?
                          1
                        :
                          2
          :
            3
      :
         (X1[7:6] <= 0)?
           (X0[7:6] <= 0)?
            3
          :
             (X1[7:5] <= 1)?
               (X1[7:4] <= 9)?
                 (X1[7:6] <= 0)?
                   (X3[7:6] <= 0)?
                    1
                  :
                     (X1[7:6] <= 0)?
                       (X3[7:6] <= 0)?
                        2
                      :
                        1
                    :
                       (X3[7:5] <= 3)?
                        2
                      :
                        1
                :
                  1
              :
                6
            :
               (X4[7:5] <= 1)?
                1
              :
                 (X3[7:6] <= 0)?
                  1
                :
                   (X3[7:4] <= 3)?
                    1
                  :
                     (X2[7:6] <= 2)?
                      1
                    :
                       (X3[7:6] <= 0)?
                         (X1[7:6] <= 0)?
                          1
                        :
                          1
                      :
                        1
        :
          4
  :
     (X4[7:6] <= 2)?
       (X3[7:4] <= 0)?
         (X0[7:6] <= 0)?
           (X2[7:6] <= 0)?
            5
          :
             (X4[7:6] <= 0)?
              1
            :
              1
        :
          2
      :
         (X1[7:6] <= 0)?
           (X2[7:6] <= 1)?
            1
          :
            1
        :
           (X4[7:3] <= 11)?
             (X2[7:6] <= 0)?
              1
            :
               (X1[7:6] <= 0)?
                 (X1[7:5] <= 0)?
                  3
                :
                  1
              :
                4
          :
             (X1[7:6] <= 1)?
               (X1[7:5] <= 4)?
                 (X1[7:6] <= 0)?
                   (X1[7:6] <= 0)?
                     (X1[7:6] <= 0)?
                      5
                    :
                       (X3[7:6] <= 1)?
                        1
                      :
                        1
                  :
                    27
                :
                   (X1[7:6] <= 0)?
                     (X2[7:5] <= 4)?
                      1
                    :
                       (X1[7:6] <= 0)?
                         (X3[7:5] <= 3)?
                          1
                        :
                          1
                      :
                         (X3[7:6] <= 2)?
                          1
                        :
                          3
                  :
                     (X1[7:5] <= 0)?
                      10
                    :
                       (X1[7:5] <= 1)?
                         (X2[7:6] <= 1)?
                          1
                        :
                          1
                      :
                         (X3[7:6] <= 0)?
                           (X1[7:6] <= 0)?
                            1
                          :
                            3
                        :
                           (X1[7:6] <= 0)?
                            19
                          :
                             (X3[7:6] <= 0)?
                              15
                            :
                               (X1[7:5] <= 1)?
                                 (X1[7:6] <= 1)?
                                   (X1[7:6] <= 0)?
                                     (X3[7:6] <= 0)?
                                      1
                                    :
                                      2
                                  :
                                     (X1[7:6] <= 0)?
                                      6
                                    :
                                       (X3[7:6] <= 2)?
                                         (X1[7:5] <= 1)?
                                          2
                                        :
                                          6
                                      :
                                         (X1[7:6] <= 0)?
                                          3
                                        :
                                          1
                                :
                                   (X1[7:6] <= 1)?
                                    18
                                  :
                                     (X3[7:5] <= 5)?
                                      4
                                    :
                                      2
                              :
                                 (X2[7:5] <= 1)?
                                  1
                                :
                                  1
              :
                41
            :
               (X1[7:6] <= 1)?
                 (X2[7:6] <= 1)?
                  2
                :
                   (X1[7:6] <= 0)?
                     (X3[7:5] <= 3)?
                      3
                    :
                      1
                  :
                    1
              :
                6
    :
       (X1[7:6] <= 1)?
        1
      :
         (X3[7:5] <= 3)?
          1
        :
           (X1[7:4] <= 5)?
            1
          :
             (X1[7:6] <= 0)?
              1
            :
              1
;
endmodule
