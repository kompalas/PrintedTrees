module top(X16, out);
input [7:0] X16;
output [3:0] out;
assign out = 
   (X16[7:5] <= 0)?
    800
  :
     (X16[7:4] <= 0)?
      794
    :
       (X16[7:4] <= -2)?
        793
      :
         (X16[7:6] <= 1)?
           (X16[7:3] <= 8)?
             (X16[7:5] <= 8)?
              734
            :
              786
          :
             (X16[7:6] <= 2)?
              738
            :
              752
        :
           (X16[7:5] <= 3)?
            805
          :
             (X16[7:2] <= 64)?
              747
            :
              745
;
endmodule
