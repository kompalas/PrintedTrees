module top(X16, out);
input [7:0] X16;
output [3:0] out;
assign out = 
   (X16[7:4] <= 0)?
    800
  :
     (X16[7:5] <= 0)?
      794
    :
       (X16[7:6] <= 0)?
        793
      :
         (X16[7:6] <= 0)?
           (X16[7:3] <= 4)?
             (X16[7:5] <= 2)?
              734
            :
              786
          :
             (X16[7:6] <= 4)?
              738
            :
              752
        :
           (X16[7:5] <= 4)?
            805
          :
             (X16[7:6] <= 2)?
              747
            :
              745
;
endmodule
