module top(X0, X1, X2, X3, X4, out);
input [7:0] X0;
input [7:0] X1;
input [7:0] X2;
input [7:0] X3;
input [7:0] X4;
output [0:0] out;
assign out = 
   (X0[7:1] <= 11)?
     (X2[7:4] <= 10)?
       (X1[7:4] <= 12)?
         (X3[7:2] <= 40)?
           (X4 <= 41)?
            1
          :
             (X1[7:5] <= 2)?
              42
            :
               (X1[7:2] <= 37)?
                 (X4[7:5] <= 7)?
                  17
                :
                   (X1[7:3] <= 15)?
                     (X1[7:4] <= 5)?
                       (X1[7:3] <= 13)?
                         (X1[7:3] <= 8)?
                           (X2[7:4] <= 6)?
                            3
                          :
                            2
                        :
                          17
                      :
                         (X0[7:4] <= 0)?
                          3
                        :
                           (X3[7:4] <= 1)?
                             (X1[7:5] <= 2)?
                               (X2[7:2] <= 9)?
                                3
                              :
                                4
                            :
                               (X2[7:5] <= 2)?
                                 (X1[7:4] <= 9)?
                                  2
                                :
                                  3
                              :
                                2
                          :
                            2
                    :
                       (X1[7:3] <= 14)?
                        40
                      :
                         (X1[7:4] <= 7)?
                           (X2[7:3] <= 4)?
                             (X1[7:4] <= 7)?
                              1
                            :
                              6
                          :
                            4
                        :
                          12
                  :
                     (X2[7:3] <= 5)?
                      2
                    :
                      1
              :
                22
        :
           (X1[7:4] <= 9)?
            5
          :
             (X3[7:4] <= 14)?
               (X2[7:3] <= 5)?
                1
              :
                 (X1[7:2] <= 33)?
                   (X1[7:5] <= 6)?
                    1
                  :
                    2
                :
                   (X1[7:5] <= 3)?
                     (X1[7:2] <= 36)?
                      1
                    :
                      1
                  :
                    2
            :
              1
      :
         (X1[7:6] <= 4)?
           (X1[7:4] <= 8)?
             (X2[7:4] <= 3)?
               (X4[7:5] <= 3)?
                1
              :
                 (X3[7:4] <= 7)?
                   (X3[7:5] <= 1)?
                     (X1[7:3] <= 21)?
                       (X1[7:1] <= 83)?
                        1
                      :
                         (X0[7:4] <= 0)?
                          1
                        :
                           (X1[7:5] <= 5)?
                            1
                          :
                            2
                    :
                      1
                  :
                    1
                :
                  1
            :
               (X3[7:3] <= 21)?
                5
              :
                1
          :
            2
        :
           (X4[7:2] <= 10)?
             (X1[7:2] <= 49)?
              1
            :
              1
          :
            9
    :
       (X1[7:5] <= 5)?
         (X1[7:3] <= 15)?
           (X1[7:3] <= 18)?
             (X1[7:5] <= 1)?
              2
            :
               (X1[7:4] <= 2)?
                1
              :
                 (X1[7:4] <= 6)?
                   (X1[7:3] <= 13)?
                     (X1[7:3] <= 9)?
                       (X3[7:4] <= 14)?
                        6
                      :
                        1
                    :
                       (X0[7:5] <= 1)?
                        1
                      :
                         (X3[7:3] <= 30)?
                           (X1[7:4] <= 10)?
                             (X3[7:5] <= 5)?
                               (X3[7:3] <= 8)?
                                 (X1[7:5] <= 3)?
                                  2
                                :
                                  2
                              :
                                 (X1[7:4] <= 5)?
                                  2
                                :
                                  1
                            :
                               (X1[7:3] <= 11)?
                                 (X4[7:3] <= 14)?
                                  1
                                :
                                  1
                              :
                                3
                          :
                            2
                        :
                          1
                  :
                     (X3[7:3] <= 29)?
                      6
                    :
                      1
                :
                   (X2[7:3] <= 27)?
                    1
                  :
                    2
          :
            6
        :
           (X1[7:4] <= 11)?
             (X1[7:4] <= 9)?
               (X4[7:3] <= 28)?
                 (X1[7:3] <= 14)?
                  1
                :
                   (X2[7:4] <= 11)?
                    1
                  :
                     (X3[7:4] <= 11)?
                      1
                    :
                      1
              :
                1
            :
               (X1[7:3] <= 17)?
                 (X3[7:5] <= 2)?
                  3
                :
                   (X1[7:5] <= 8)?
                    1
                  :
                     (X3[7:5] <= 7)?
                       (X2[7:4] <= 13)?
                        1
                      :
                        1
                    :
                      2
              :
                 (X3[7:4] <= 5)?
                  1
                :
                   (X4[7:1] <= 68)?
                    1
                  :
                     (X0[7:1] <= 8)?
                      1
                    :
                       (X3[7:1] <= 112)?
                         (X1[7:3] <= 21)?
                           (X3[7:3] <= 22)?
                            2
                          :
                             (X1[7:4] <= 9)?
                               (X2[7:2] <= 52)?
                                1
                              :
                                1
                            :
                              2
                        :
                           (X2[7:4] <= 13)?
                            2
                          :
                             (X1[7:3] <= 17)?
                               (X3[7:4] <= 10)?
                                1
                              :
                                1
                            :
                              1
                      :
                         (X1[7:5] <= 5)?
                          1
                        :
                          2
          :
            3
      :
         (X1[7:4] <= 11)?
           (X0[7:3] <= 6)?
            3
          :
             (X1[7:4] <= 13)?
               (X1[7:3] <= 22)?
                 (X1[7:3] <= 19)?
                   (X3[7:3] <= 13)?
                    1
                  :
                     (X1[7:5] <= 4)?
                       (X3 <= 223)?
                        2
                      :
                        1
                    :
                       (X3 <= 229)?
                        2
                      :
                        1
                :
                  1
              :
                6
            :
               (X4[7:4] <= 8)?
                1
              :
                 (X3[7:1] <= 17)?
                  1
                :
                   (X3[7:4] <= 4)?
                    1
                  :
                     (X2[7:2] <= 54)?
                      1
                    :
                       (X3[7:4] <= 11)?
                         (X1[7:3] <= 22)?
                          1
                        :
                          1
                      :
                        1
        :
          4
  :
     (X4[7:1] <= 105)?
       (X3[7:4] <= 1)?
         (X0[7:6] <= 4)?
           (X2[7:4] <= 9)?
            5
          :
             (X4[7:4] <= 6)?
              1
            :
              1
        :
          2
      :
         (X1[7:3] <= 5)?
           (X2[7:4] <= 11)?
            1
          :
            1
        :
           (X4[7:3] <= 21)?
             (X2[7:4] <= 9)?
              1
            :
               (X1[7:1] <= 70)?
                 (X1[7:5] <= 5)?
                  3
                :
                  1
              :
                4
          :
             (X1[7:4] <= 14)?
               (X1[7:2] <= 44)?
                 (X1[7:3] <= 16)?
                   (X1[7:3] <= 10)?
                     (X1[7:2] <= 16)?
                      5
                    :
                       (X3[7:4] <= 14)?
                        1
                      :
                        1
                  :
                    27
                :
                   (X1[7:1] <= 60)?
                     (X2[7:3] <= 28)?
                      1
                    :
                       (X1[7:4] <= 6)?
                         (X3[7:3] <= 27)?
                          1
                        :
                          1
                      :
                         (X3 <= 162)?
                          1
                        :
                          3
                  :
                     (X1[7:4] <= 10)?
                      10
                    :
                       (X1[7:4] <= 9)?
                         (X2[7:1] <= 87)?
                          1
                        :
                          1
                      :
                         (X3[7:3] <= 12)?
                           (X1[7:4] <= 7)?
                            1
                          :
                            3
                        :
                           (X1[7:4] <= 9)?
                            19
                          :
                             (X3[7:5] <= 4)?
                              15
                            :
                               (X1[7:2] <= 44)?
                                 (X1[7:4] <= 12)?
                                   (X1[7:4] <= 10)?
                                     (X3[7:3] <= 28)?
                                      1
                                    :
                                      2
                                  :
                                     (X1[7:3] <= 21)?
                                      6
                                    :
                                       (X3[7:4] <= 14)?
                                         (X1[7:4] <= 10)?
                                          2
                                        :
                                          6
                                      :
                                         (X1[7:4] <= 10)?
                                          3
                                        :
                                          1
                                :
                                   (X1[7:4] <= 11)?
                                    18
                                  :
                                     (X3[7:3] <= 28)?
                                      4
                                    :
                                      2
                              :
                                 (X2[7:1] <= 85)?
                                  1
                                :
                                  1
              :
                41
            :
               (X1[7:1] <= 112)?
                 (X2[7:5] <= 6)?
                  2
                :
                   (X1[7:4] <= 16)?
                     (X3[7:4] <= 15)?
                      3
                    :
                      1
                  :
                    1
              :
                6
    :
       (X1[7:2] <= 30)?
        1
      :
         (X3[7:5] <= 5)?
          1
        :
           (X1[7:5] <= 4)?
            1
          :
             (X1[7:5] <= 3)?
              1
            :
              1
;
endmodule
