module top(X0, X1, X2, X3, X4, X5, X6, X7, X8, out);
input [7:0] X0;
input [7:0] X1;
input [7:0] X2;
input [7:0] X3;
input [7:0] X4;
input [7:0] X5;
input [7:0] X6;
input [7:0] X7;
input [7:0] X8;
output [1:0] out;
assign out = 
   (X2 <= 71)?
     (X6 <= 43)?
       (X5 <= 100)?
        291
      :
         (X3 <= 43)?
          2
        :
          2
    :
       (X7 <= 14)?
        10
      :
         (X1 <= 156)?
           (X5 <= 100)?
             (X3 <= 100)?
               (X0 <= 19)?
                5
              :
                 (X6 <= 71)?
                  3
                :
                   (X4 <= 171)?
                    3
                  :
                    1
            :
              2
          :
            5
        :
          9
  :
     (X7 <= 100)?
       (X6 <= 213)?
         (X1 <= 213)?
           (X4 <= 128)?
             (X8 <= 185)?
               (X3 <= 228)?
                 (X5 <= 128)?
                  5
                :
                   (X6 <= 128)?
                    1
                  :
                    1
              :
                1
            :
              3
          :
            5
        :
          7
      :
        21
    :
      101
;
endmodule
