module top(X0, X1, X2, X3, X4, X5, X6, X7, X8, X9, X10, out);
input [7:0] X0;
input [7:0] X1;
input [7:0] X2;
input [7:0] X3;
input [7:0] X4;
input [7:0] X5;
input [7:0] X6;
input [7:0] X7;
input [7:0] X8;
input [7:0] X9;
input [7:0] X10;
output [3:0] out;
assign out = 
   (X10[7:6] <= 1)?
     (X9[7:6] <= 0)?
       (X6[7:6] <= 0)?
         (X1[7:6] <= 0)?
           (X9[7:6] <= 0)?
            16
          :
             (X7[7:6] <= 1)?
               (X10[7:5] <= 0)?
                1
              :
                7
            :
               (X5[7:6] <= 0)?
                 (X5[7:6] <= 0)?
                   (X10[7:6] <= 0)?
                    10
                  :
                     (X10[7:4] <= 1)?
                       (X7[7:6] <= 0)?
                         (X4[7:6] <= 0)?
                          1
                        :
                          4
                      :
                        1
                    :
                      3
                :
                   (X1[7:6] <= 0)?
                    1
                  :
                     (X7[7:6] <= 1)?
                      2
                    :
                       (X6[7:6] <= 0)?
                         (X1[7:5] <= 0)?
                           (X6[7:5] <= 0)?
                            1
                          :
                            1
                        :
                          11
                      :
                         (X1[7:6] <= 0)?
                          3
                        :
                           (X3[7:6] <= 0)?
                             (X1[7:6] <= 0)?
                              1
                            :
                              2
                          :
                            3
              :
                 (X4[7:6] <= 0)?
                   (X5[7:6] <= 0)?
                    1
                  :
                    2
                :
                  3
        :
           (X0[7:6] <= 0)?
             (X1[7:5] <= 1)?
               (X2[7:6] <= 0)?
                3
              :
                 (X4[7:6] <= 0)?
                  4
                :
                  2
            :
               (X7[7:6] <= 0)?
                 (X4[7:6] <= 3)?
                  1
                :
                  1
              :
                 (X10[7:6] <= 0)?
                   (X6[7:6] <= 0)?
                    26
                  :
                    1
                :
                  1
          :
             (X6[7:6] <= 0)?
               (X9[7:6] <= 0)?
                 (X1[7:4] <= 3)?
                  7
                :
                   (X7[7:6] <= 0)?
                    1
                  :
                    5
              :
                 (X7[7:6] <= 0)?
                   (X7[7:5] <= 1)?
                     (X6[7:6] <= 0)?
                       (X7[7:6] <= 0)?
                        2
                      :
                        1
                    :
                      4
                  :
                    3
                :
                  12
            :
               (X2[7:5] <= 1)?
                3
              :
                 (X3[7:5] <= 1)?
                  2
                :
                   (X8[7:6] <= 1)?
                    1
                  :
                    1
      :
         (X10[7:6] <= 0)?
           (X5[7:6] <= 0)?
             (X3[7:5] <= 0)?
               (X8[7:6] <= 0)?
                1
              :
                1
            :
              13
          :
             (X3[7:6] <= 0)?
               (X6[7:6] <= 0)?
                 (X8[7:6] <= 4)?
                   (X2[7:6] <= 0)?
                    17
                  :
                     (X2[7:6] <= 0)?
                       (X8[7:6] <= 1)?
                        7
                      :
                         (X9[7:6] <= 0)?
                           (X8[7:6] <= 0)?
                             (X7[7:6] <= 0)?
                               (X1[7:5] <= 1)?
                                1
                              :
                                4
                            :
                              5
                          :
                             (X0[7:6] <= 0)?
                               (X0[7:6] <= 0)?
                                3
                              :
                                2
                            :
                              14
                        :
                          3
                    :
                       (X1[7:6] <= 0)?
                        1
                      :
                        20
                :
                  2
              :
                26
            :
              2
        :
           (X6[7:6] <= 0)?
            2
          :
             (X3[7:6] <= 0)?
              1
            :
              1
    :
       (X6[7:6] <= 0)?
         (X1[7:6] <= 0)?
           (X10[7:5] <= 0)?
             (X0[7:6] <= 0)?
               (X2[7:6] <= 0)?
                 (X8[7:6] <= 2)?
                   (X7[7:6] <= 0)?
                    2
                  :
                     (X4[7:6] <= 0)?
                       (X9[7:6] <= 0)?
                         (X8[7:6] <= 0)?
                          1
                        :
                          1
                      :
                        17
                    :
                       (X0[7:6] <= 0)?
                        2
                      :
                        3
                :
                  3
              :
                7
            :
              11
          :
             (X9[7:6] <= 0)?
               (X8[7:4] <= 2)?
                 (X7[7:6] <= 0)?
                  3
                :
                  2
              :
                 (X2[7:6] <= 0)?
                   (X0[7:5] <= 0)?
                     (X7[7:6] <= 0)?
                      1
                    :
                      5
                  :
                     (X4[7:6] <= 0)?
                       (X8[7:6] <= 0)?
                        1
                      :
                        7
                    :
                      2
                :
                   (X2[7:6] <= 0)?
                    8
                  :
                     (X5[7:6] <= 0)?
                       (X5[7:6] <= 0)?
                        2
                      :
                         (X10[7:5] <= 0)?
                          1
                        :
                          3
                    :
                      4
            :
               (X5[7:5] <= 0)?
                 (X4[7:6] <= 0)?
                  2
                :
                  3
              :
                 (X5[7:6] <= 0)?
                   (X4[7:6] <= 0)?
                     (X7[7:6] <= 2)?
                      1
                    :
                      3
                  :
                    2
                :
                  8
        :
           (X8[7:4] <= 7)?
             (X0[7:6] <= 0)?
               (X8[7:6] <= 1)?
                 (X10[7:6] <= 0)?
                   (X9[7:4] <= 8)?
                     (X2[7:4] <= 3)?
                      23
                    :
                       (X9[7:6] <= 0)?
                         (X0[7:6] <= 0)?
                          3
                        :
                          1
                      :
                         (X8[7:6] <= 0)?
                          1
                        :
                          12
                  :
                     (X1[7:5] <= 0)?
                      1
                    :
                      1
                :
                   (X9[7:6] <= 0)?
                     (X1[7:6] <= 0)?
                       (X10[7:6] <= 0)?
                        2
                      :
                        5
                    :
                      8
                  :
                    7
              :
                 (X1[7:6] <= 0)?
                   (X2[7:6] <= 0)?
                     (X10[7:6] <= 0)?
                      8
                    :
                       (X9[7:6] <= 0)?
                         (X8[7:5] <= 3)?
                           (X3[7:5] <= 0)?
                             (X10[7:5] <= 0)?
                               (X6[7:5] <= 0)?
                                 (X3[7:6] <= 0)?
                                   (X8[7:6] <= 2)?
                                     (X5[7:6] <= 0)?
                                       (X5[7:6] <= 0)?
                                         (X5[7:6] <= 0)?
                                          2
                                        :
                                           (X9[7:4] <= 0)?
                                            5
                                          :
                                            1
                                      :
                                         (X0[7:6] <= 0)?
                                          3
                                        :
                                          1
                                    :
                                      3
                                  :
                                    6
                                :
                                   (X1[7:6] <= 0)?
                                    12
                                  :
                                    4
                              :
                                10
                            :
                               (X6[7:6] <= 0)?
                                 (X8[7:6] <= 0)?
                                  5
                                :
                                   (X2[7:6] <= 0)?
                                    3
                                  :
                                     (X1[7:6] <= 0)?
                                      2
                                    :
                                       (X7[7:6] <= 0)?
                                         (X4[7:6] <= 0)?
                                          7
                                        :
                                          1
                                      :
                                         (X6[7:6] <= 0)?
                                          1
                                        :
                                          2
                              :
                                9
                          :
                            6
                        :
                           (X6[7:6] <= 0)?
                             (X7[7:6] <= 0)?
                              1
                            :
                               (X5[7:6] <= 0)?
                                2
                              :
                                1
                          :
                            7
                      :
                        8
                  :
                     (X5[7:6] <= 0)?
                      7
                    :
                      1
                :
                   (X3[7:6] <= 0)?
                    1
                  :
                    1
            :
               (X4[7:6] <= 0)?
                 (X8[7:6] <= 0)?
                   (X2[7:6] <= 0)?
                     (X3[7:6] <= 0)?
                       (X10[7:6] <= 0)?
                        2
                      :
                        1
                    :
                      2
                  :
                     (X9[7:6] <= 0)?
                      3
                    :
                      1
                :
                   (X5[7:6] <= 0)?
                    3
                  :
                     (X8[7:6] <= 0)?
                      8
                    :
                       (X9[7:6] <= 0)?
                        1
                      :
                         (X5[7:4] <= 2)?
                          6
                        :
                           (X7[7:6] <= 0)?
                            1
                          :
                            1
              :
                 (X5[7:6] <= 0)?
                  2
                :
                  1
          :
             (X5[7:6] <= 0)?
               (X7[7:6] <= 0)?
                 (X9[7:6] <= 0)?
                  2
                :
                  1
              :
                 (X9[7:6] <= 0)?
                  1
                :
                  2
            :
               (X3[7:6] <= 0)?
                16
              :
                1
      :
         (X9[7:6] <= 1)?
           (X3[7:5] <= 2)?
             (X1[7:5] <= 0)?
              1
            :
               (X9[7:6] <= 0)?
                 (X5[7:5] <= 1)?
                  2
                :
                  7
              :
                 (X3[7:5] <= 0)?
                  1
                :
                   (X6[7:6] <= 0)?
                     (X4[7:5] <= 0)?
                      1
                    :
                      3
                  :
                    48
          :
            2
        :
           (X10[7:6] <= 0)?
            2
          :
            4
  :
     (X9[7:6] <= 0)?
       (X1[7:6] <= 0)?
         (X1[7:6] <= 0)?
           (X8[7:5] <= 0)?
             (X7[7:3] <= 13)?
               (X3[7:5] <= 0)?
                 (X2[7:6] <= 0)?
                   (X6[7:5] <= 0)?
                    5
                  :
                     (X2[7:6] <= 0)?
                       (X10[7:6] <= 0)?
                        2
                      :
                        1
                    :
                      5
                :
                   (X10[7:5] <= 1)?
                     (X8[7:6] <= 0)?
                      1
                    :
                      1
                  :
                    9
              :
                5
            :
               (X4[7:6] <= 0)?
                3
              :
                3
          :
             (X7[7:5] <= 0)?
               (X7[7:6] <= 0)?
                 (X7[7:6] <= 0)?
                  3
                :
                  2
              :
                16
            :
               (X4[7:6] <= 0)?
                 (X10[7:6] <= 0)?
                  3
                :
                  2
              :
                 (X4[7:6] <= 0)?
                   (X8[7:5] <= 3)?
                    2
                  :
                    2
                :
                  5
        :
           (X5[7:6] <= 0)?
             (X3[7:6] <= 0)?
               (X7[7:5] <= 2)?
                 (X1[7:6] <= 0)?
                  1
                :
                   (X6[7:6] <= 0)?
                    3
                  :
                     (X1[7:6] <= 0)?
                       (X7[7:5] <= 1)?
                        1
                      :
                        7
                    :
                      2
              :
                 (X2[7:6] <= 0)?
                  2
                :
                  1
            :
              10
          :
             (X6[7:6] <= 0)?
               (X10[7:6] <= 0)?
                 (X7[7:6] <= 0)?
                  4
                :
                  1
              :
                4
            :
               (X9[7:6] <= 1)?
                 (X3[7:6] <= 0)?
                   (X5[7:6] <= 0)?
                    7
                  :
                     (X7[7:5] <= 0)?
                       (X6[7:6] <= 0)?
                        3
                      :
                        1
                    :
                       (X5[7:6] <= 0)?
                        4
                      :
                         (X10[7:6] <= 0)?
                          1
                        :
                          1
                :
                   (X1[7:6] <= 0)?
                    3
                  :
                    1
              :
                 (X5[7:6] <= 0)?
                   (X4[7:6] <= 0)?
                     (X7[7:6] <= 0)?
                      2
                    :
                      3
                  :
                     (X2[7:6] <= 0)?
                      24
                    :
                       (X7[7:6] <= 0)?
                        1
                      :
                        1
                :
                  2
      :
         (X3[7:6] <= 0)?
          2
        :
           (X9[7:5] <= 0)?
            3
          :
            3
    :
       (X10[7:6] <= 0)?
         (X1[7:5] <= 0)?
           (X6[7:6] <= 0)?
             (X8[7:4] <= 5)?
               (X0[7:5] <= 0)?
                 (X1[7:6] <= 0)?
                   (X8[7:4] <= 3)?
                    4
                  :
                    1
                :
                   (X2[7:5] <= 3)?
                    1
                  :
                    2
              :
                 (X1[7:6] <= 0)?
                  11
                :
                  1
            :
               (X6[7:6] <= 0)?
                 (X3[7:6] <= 0)?
                   (X9[7:6] <= 1)?
                    3
                  :
                    2
                :
                  3
              :
                 (X9[7:6] <= 1)?
                  6
                :
                   (X8[7:6] <= 4)?
                     (X8[7:6] <= 0)?
                       (X1[7:6] <= 0)?
                        1
                      :
                        2
                    :
                      5
                  :
                    5
          :
             (X0[7:5] <= 2)?
               (X4[7:6] <= 0)?
                 (X9[7:6] <= 0)?
                  2
                :
                  1
              :
                6
            :
               (X2[7:6] <= 0)?
                3
              :
                1
        :
           (X4[7:6] <= 0)?
             (X3[7:6] <= 0)?
               (X1[7:5] <= 0)?
                 (X8[7:6] <= 0)?
                   (X3[7:6] <= 0)?
                     (X6[7:6] <= 0)?
                      1
                    :
                      6
                  :
                    1
                :
                  28
              :
                 (X1[7:6] <= 0)?
                  3
                :
                  7
            :
               (X8[7:6] <= 0)?
                 (X9[7:5] <= 0)?
                  10
                :
                   (X9[7:5] <= 2)?
                    2
                  :
                    1
              :
                 (X7[7:5] <= 0)?
                   (X10[7:6] <= 0)?
                    3
                  :
                     (X1[7:5] <= 0)?
                      1
                    :
                      1
                :
                  5
          :
             (X0[7:4] <= 3)?
               (X3[7:6] <= 0)?
                3
              :
                1
            :
               (X6[7:6] <= 0)?
                7
              :
                 (X0[7:5] <= 1)?
                  2
                :
                  2
      :
         (X6[7:6] <= 0)?
           (X4[7:6] <= 0)?
             (X4[7:6] <= 0)?
               (X1[7:6] <= 0)?
                7
              :
                 (X9[7:4] <= 0)?
                  1
                :
                  4
            :
               (X6[7:6] <= 0)?
                 (X9[7:6] <= 0)?
                  1
                :
                  5
              :
                 (X1[7:6] <= 0)?
                  3
                :
                  1
          :
            10
        :
           (X9[7:4] <= 2)?
             (X8[7:6] <= 1)?
               (X5[7:5] <= 0)?
                15
              :
                1
            :
               (X4[7:6] <= 0)?
                 (X4[7:6] <= 0)?
                  2
                :
                   (X6[7:6] <= 0)?
                    1
                  :
                    2
              :
                 (X10[7:5] <= 3)?
                  1
                :
                  2
          :
             (X5[7:6] <= 0)?
               (X8[7:6] <= 2)?
                 (X7[7:6] <= 0)?
                  2
                :
                   (X10[7:5] <= 2)?
                    2
                  :
                    1
              :
                 (X1[7:6] <= 2)?
                   (X7[7:6] <= 0)?
                    20
                  :
                     (X8[7:6] <= 2)?
                      2
                    :
                      1
                :
                  1
            :
               (X8[7:6] <= 0)?
                 (X10[7:6] <= 1)?
                   (X4[7:6] <= 0)?
                    5
                  :
                     (X7[7:6] <= 0)?
                      5
                    :
                      4
                :
                  1
              :
                 (X6[7:5] <= 0)?
                   (X1[7:6] <= 0)?
                    2
                  :
                    1
                :
                  8
;
endmodule
