module top(X2, X6, X9, X10, X12, X14, X23, X28, X32, X36, X37, X40, X41, X42, X43, X50, X51, X54, X55, X56, X57, X58, X63, X65, X68, X69, X74, X76, X77, X86, X88, X89, X100, X102, X111, X115, X117, X118, X128, X131, X133, X139, X140, X141, X144, X145, X147, X150, X152, X158, X175, X178, X179, X181, X185, X187, X189, X196, X197, X198, X203, X204, X214, X221, X224, X230, X238, X243, X246, X252, X257, X264, X266, X270, X276, X280, X288, X293, X295, X300, X301, X302, X305, X306, X317, X321, X330, X331, X335, X339, X343, X357, X358, X365, X369, X371, X374, X387, X390, X394, X396, X407, X410, X415, X417, X418, X427, X434, X435, X440, X448, X449, X453, X454, X464, X467, X476, X485, X486, X490, X491, X492, X494, X498, X504, X507, X509, X510, X515, X536, X546, X552, X554, X555, X557, X558, X559, X560, out);
input [7:0] X2;
input [7:0] X6;
input [7:0] X9;
input [7:0] X10;
input [7:0] X12;
input [7:0] X14;
input [7:0] X23;
input [7:0] X28;
input [7:0] X32;
input [7:0] X36;
input [7:0] X37;
input [7:0] X40;
input [7:0] X41;
input [7:0] X42;
input [7:0] X43;
input [7:0] X50;
input [7:0] X51;
input [7:0] X54;
input [7:0] X55;
input [7:0] X56;
input [7:0] X57;
input [7:0] X58;
input [7:0] X63;
input [7:0] X65;
input [7:0] X68;
input [7:0] X69;
input [7:0] X74;
input [7:0] X76;
input [7:0] X77;
input [7:0] X86;
input [7:0] X88;
input [7:0] X89;
input [7:0] X100;
input [7:0] X102;
input [7:0] X111;
input [7:0] X115;
input [7:0] X117;
input [7:0] X118;
input [7:0] X128;
input [7:0] X131;
input [7:0] X133;
input [7:0] X139;
input [7:0] X140;
input [7:0] X141;
input [7:0] X144;
input [7:0] X145;
input [7:0] X147;
input [7:0] X150;
input [7:0] X152;
input [7:0] X158;
input [7:0] X175;
input [7:0] X178;
input [7:0] X179;
input [7:0] X181;
input [7:0] X185;
input [7:0] X187;
input [7:0] X189;
input [7:0] X196;
input [7:0] X197;
input [7:0] X198;
input [7:0] X203;
input [7:0] X204;
input [7:0] X214;
input [7:0] X221;
input [7:0] X224;
input [7:0] X230;
input [7:0] X238;
input [7:0] X243;
input [7:0] X246;
input [7:0] X252;
input [7:0] X257;
input [7:0] X264;
input [7:0] X266;
input [7:0] X270;
input [7:0] X276;
input [7:0] X280;
input [7:0] X288;
input [7:0] X293;
input [7:0] X295;
input [7:0] X300;
input [7:0] X301;
input [7:0] X302;
input [7:0] X305;
input [7:0] X306;
input [7:0] X317;
input [7:0] X321;
input [7:0] X330;
input [7:0] X331;
input [7:0] X335;
input [7:0] X339;
input [7:0] X343;
input [7:0] X357;
input [7:0] X358;
input [7:0] X365;
input [7:0] X369;
input [7:0] X371;
input [7:0] X374;
input [7:0] X387;
input [7:0] X390;
input [7:0] X394;
input [7:0] X396;
input [7:0] X407;
input [7:0] X410;
input [7:0] X415;
input [7:0] X417;
input [7:0] X418;
input [7:0] X427;
input [7:0] X434;
input [7:0] X435;
input [7:0] X440;
input [7:0] X448;
input [7:0] X449;
input [7:0] X453;
input [7:0] X454;
input [7:0] X464;
input [7:0] X467;
input [7:0] X476;
input [7:0] X485;
input [7:0] X486;
input [7:0] X490;
input [7:0] X491;
input [7:0] X492;
input [7:0] X494;
input [7:0] X498;
input [7:0] X504;
input [7:0] X507;
input [7:0] X509;
input [7:0] X510;
input [7:0] X515;
input [7:0] X536;
input [7:0] X546;
input [7:0] X552;
input [7:0] X554;
input [7:0] X555;
input [7:0] X557;
input [7:0] X558;
input [7:0] X559;
input [7:0] X560;
output [2:0] out;
assign out = 
   (X102[7:3] <= 20)?
     (X56[7:2] <= 18)?
       (X63[7:3] <= 8)?
         (X118[7:3] <= 27)?
           (X88[7:3] <= 12)?
            336
          :
            1
        :
           (X293[7:4] <= 9)?
            3
          :
            3
      :
         (X54[7:3] <= 27)?
           (X51[7:2] <= 49)?
            16
          :
             (X198[7:5] <= 3)?
              4
            :
              24
        :
           (X55[7:4] <= 9)?
            7
          :
            25
    :
       (X51[7:2] <= 33)?
         (X139 <= 1)?
           (X58[7:2] <= 3)?
             (X139[7:2] <= 0)?
              53
            :
               (X417[7:3] <= 1)?
                 (X57[7:4] <= 1)?
                   (X453[7:3] <= 17)?
                    28
                  :
                     (X252[7:2] <= 0)?
                      8
                    :
                      3
                :
                   (X306[7:4] <= 1)?
                    15
                  :
                    2
              :
                 (X14[7:4] <= 16)?
                   (X305[7:3] <= 0)?
                    3
                  :
                    2
                :
                  54
          :
             (X41[7:4] <= 6)?
              14
            :
              29
        :
           (X181[7:3] <= 2)?
             (X51[7:3] <= 13)?
               (X54[7:2] <= 9)?
                11
              :
                 (X50[7:3] <= 17)?
                   (X448[7:3] <= 7)?
                     (X435[7:4] <= 2)?
                       (X147[7:5] <= 7)?
                         (X536[7:4] <= 11)?
                          32
                        :
                          1
                      :
                         (X554[7:3] <= 17)?
                          6
                        :
                          3
                    :
                       (X115[7:4] <= 7)?
                         (X144[7:3] <= 14)?
                           (X357[7:2] <= 3)?
                            3
                          :
                            4
                        :
                          26
                      :
                        256
                  :
                     (X115[7:4] <= 7)?
                       (X485[7:3] <= 0)?
                        8
                      :
                        2
                    :
                      8
                :
                   (X559[7:3] <= 15)?
                     (X187[7:3] <= 8)?
                      1
                    :
                      37
                  :
                     (X54[7:2] <= 21)?
                       (X23[7:3] <= 6)?
                        2
                      :
                        8
                    :
                       (X434[7:4] <= 3)?
                        24
                      :
                        1
            :
               (X560[7:4] <= 10)?
                 (X40[7:3] <= 32)?
                   (X32[7:4] <= 11)?
                    45
                  :
                     (X14[7:3] <= 30)?
                       (X557[7:3] <= 5)?
                        1
                      :
                        4
                    :
                      8
                :
                  10
              :
                 (X189[7:4] <= 6)?
                   (X492[7:2] <= 0)?
                    1
                  :
                    35
                :
                   (X224[7:4] <= 7)?
                    6
                  :
                     (X300[7:5] <= 4)?
                       (X554[7:3] <= 25)?
                        3
                      :
                        1
                    :
                      13
          :
             (X150[7:3] <= 20)?
               (X498[7:3] <= 0)?
                3
              :
                4
            :
               (X196[7:3] <= 15)?
                 (X214[7:4] <= 8)?
                  3
                :
                  1
              :
                6
      :
         (X57[7:3] <= 0)?
           (X41[7:5] <= 3)?
            18
          :
             (X145[7:2] <= 37)?
               (X41[7:3] <= 15)?
                7
              :
                8
            :
              54
        :
           (X179[7:2] <= 6)?
             (X36[7:3] <= 7)?
               (X214[7:4] <= 1)?
                3
              :
                2
            :
              232
          :
             (X427[7:4] <= 3)?
              2
            :
              3
  :
     (X65[7:4] <= 5)?
       (X69[7:4] <= 6)?
         (X560[7:3] <= 17)?
           (X371[7:3] <= 13)?
             (X264[7:3] <= 13)?
              2
            :
              5
          :
             (X494[7:3] <= 1)?
              10
            :
               (X65[7:4] <= 2)?
                2
              :
                2
        :
           (X330[7:3] <= 1)?
             (X490[7:5] <= 1)?
              18
            :
               (X507[7:2] <= 13)?
                1
              :
                3
          :
             (X158[7:2] <= 38)?
               (X246[7:3] <= 12)?
                 (X515[7:4] <= 10)?
                  109
                :
                  1
              :
                 (X203[7:4] <= 7)?
                  2
                :
                   (X407[7:3] <= 4)?
                    1
                  :
                    1
            :
               (X486[7:2] <= 4)?
                 (X12[7:2] <= 47)?
                   (X89[7:3] <= 10)?
                     (X491[7:4] <= 2)?
                      12
                    :
                      1
                  :
                     (X302[7:3] <= 11)?
                      10
                    :
                      1
                :
                   (X331[7:3] <= 2)?
                    1
                  :
                    4
              :
                25
      :
         (X330[7:3] <= 1)?
           (X434[7:4] <= 3)?
             (X28[7:3] <= 15)?
               (X343[7:4] <= 3)?
                2
              :
                 (X270[7:2] <= 11)?
                  2
                :
                  2
            :
               (X77[7:2] <= 64)?
                103
              :
                1
          :
             (X276[7:3] <= 3)?
              7
            :
               (X185[7:3] <= 24)?
                10
              :
                1
        :
           (X57[7:3] <= 1)?
             (X257[7:2] <= 44)?
               (X464[7:3] <= 1)?
                 (X175[7:2] <= 20)?
                   (X74[7:2] <= 51)?
                    4
                  :
                    2
                :
                   (X288[7:4] <= 14)?
                    8
                  :
                    1
              :
                 (X390[7:3] <= 2)?
                  1
                :
                  31
            :
               (X335[7:2] <= 5)?
                2
              :
                21
          :
             (X14[7:2] <= 29)?
               (X374[7:2] <= 16)?
                5
              :
                34
            :
               (X40[7:4] <= 16)?
                 (X76[7:3] <= 24)?
                  3
                :
                   (X140[7:3] <= 9)?
                    14
                  :
                    2
              :
                 (X203[7:3] <= 8)?
                   (X41[7:3] <= 20)?
                    3
                  :
                    10
                :
                   (X552[7:3] <= 18)?
                     (X238[7:5] <= 6)?
                       (X295[7:4] <= 4)?
                         (X141[7:3] <= 5)?
                          1
                        :
                          20
                      :
                         (X230[7:2] <= 17)?
                           (X117[7:4] <= 5)?
                            1
                          :
                            8
                        :
                          6
                    :
                       (X56[7:2] <= 59)?
                        72
                      :
                        1
                  :
                     (X243[7:4] <= 3)?
                      1
                    :
                      4
    :
       (X509[7:2] <= 23)?
         (X37[7:2] <= 42)?
           (X476[7:3] <= 0)?
             (X394[7:4] <= 2)?
               (X102[7:4] <= 15)?
                 (X560[7:4] <= 12)?
                  3
                :
                   (X221[7:3] <= 26)?
                     (X339[7:3] <= 2)?
                      4
                    :
                      4
                  :
                    57
              :
                3
            :
               (X317[7:3] <= 3)?
                 (X449[7:3] <= 4)?
                   (X387[7:1] <= 1)?
                    2
                  :
                    39
                :
                   (X102[7:4] <= 15)?
                    8
                  :
                     (X396[7:3] <= 2)?
                      1
                    :
                      2
              :
                 (X427[7:4] <= 4)?
                   (X100[7:3] <= 11)?
                    24
                  :
                     (X369[7:5] <= 2)?
                       (X152[7:3] <= 18)?
                        2
                      :
                        7
                    :
                      13
                :
                   (X178[7:3] <= 1)?
                     (X358[7:3] <= 1)?
                      1
                    :
                      8
                  :
                     (X204[7:4] <= 1)?
                       (X266[7:2] <= 28)?
                        3
                      :
                        1
                    :
                       (X128[7:3] <= 5)?
                         (X546[7:3] <= 7)?
                          1
                        :
                          2
                      :
                        17
          :
             (X41[7:2] <= 20)?
              13
            :
               (X42[7:3] <= 17)?
                 (X559[7:3] <= 15)?
                   (X43[7:3] <= 2)?
                     (X440[7:3] <= 4)?
                       (X10[7:4] <= 4)?
                         (X510[7:4] <= 13)?
                          4
                        :
                          3
                      :
                        69
                    :
                      3
                  :
                     (X28[7:2] <= 41)?
                       (X68[7:4] <= 13)?
                         (X418[7:2] <= 14)?
                          11
                        :
                          2
                      :
                        4
                    :
                       (X280[7:3] <= 13)?
                        3
                      :
                        7
                :
                   (X434[7:2] <= 8)?
                     (X6[7:3] <= 10)?
                       (X133[7:4] <= 13)?
                         (X558[7:5] <= 0)?
                          3
                        :
                          1
                      :
                        46
                    :
                      7
                  :
                     (X467[7:3] <= 1)?
                       (X68[7:4] <= 14)?
                        4
                      :
                        2
                    :
                       (X555[7:3] <= 3)?
                         (X2[7:3] <= 10)?
                          2
                        :
                          9
                      :
                        192
              :
                 (X111[7:2] <= 39)?
                  5
                :
                  5
        :
           (X55[7:3] <= 23)?
             (X197[7:3] <= 15)?
               (X41[7:3] <= 15)?
                 (X415[7:2] <= 3)?
                  1
                :
                  1
              :
                23
            :
               (X2[7:5] <= 3)?
                4
              :
                 (X50[7:3] <= 21)?
                  20
                :
                   (X86[7:3] <= 13)?
                    1
                  :
                    1
          :
             (X41[7:4] <= 10)?
               (X158[7:3] <= 25)?
                27
              :
                 (X454[7:3] <= 15)?
                  1
                :
                  1
            :
              17
      :
         (X9[7:3] <= 17)?
           (X50[7:2] <= 21)?
            9
          :
             (X276[7:2] <= 16)?
               (X321[7:4] <= 2)?
                 (X560[7:3] <= 27)?
                  32
                :
                  2
              :
                 (X504[7:3] <= 15)?
                   (X410[7:3] <= 7)?
                     (X365[7:4] <= 8)?
                      3
                    :
                      13
                  :
                     (X301[7:2] <= 2)?
                      1
                    :
                      5
                :
                  13
            :
               (X131[7:3] <= 3)?
                1
              :
                7
        :
          66
;
endmodule
