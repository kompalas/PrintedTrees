module top(X16, out);
input [7:0] X16;
output [3:0] out;
assign out = 
   (X16[7:6] <= 1)?
    796
  :
     (X16[7:6] <= 1)?
       (X16[7:6] <= 1)?
        785
      :
        815
    :
       (X16[7:6] <= 3)?
         (X16[7:2] <= 31)?
           (X16[7:4] <= 7)?
            711
          :
            799
        :
           (X16[7:6] <= 4)?
            749
          :
            752
      :
         (X16[7:5] <= 7)?
          831
        :
           (X16[7:3] <= 31)?
            747
          :
            709
;
endmodule
