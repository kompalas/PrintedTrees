module top(X0, X1, X2, X3, X4, X5, out);
input [7:0] X0;
input [7:0] X1;
input [7:0] X2;
input [7:0] X3;
input [7:0] X4;
input [7:0] X5;
output [1:0] out;
assign out = 
   (X5[7:2] <= 3)?
     (X3[7:5] <= 3)?
       (X4[7:1] <= 66)?
        13
      :
         (X1[7:3] <= 10)?
           (X0[7:3] <= 2)?
            1
          :
            11
        :
           (X4[7:3] <= 19)?
             (X1[7:4] <= 7)?
               (X0[7:3] <= 5)?
                 (X5[7:3] <= 1)?
                  8
                :
                   (X4[7:3] <= 21)?
                    1
                  :
                    1
              :
                 (X3[7:2] <= 14)?
                  3
                :
                   (X0[7:3] <= 7)?
                    1
                  :
                    4
            :
              6
          :
             (X5[7:2] <= 5)?
               (X1[7:3] <= 15)?
                7
              :
                1
            :
              2
    :
       (X4[7:4] <= 8)?
         (X3[7:3] <= 11)?
           (X1[7:3] <= 18)?
             (X4[7:2] <= 28)?
              6
            :
               (X5[7:4] <= 1)?
                 (X5[7:1] <= 1)?
                  1
                :
                  3
              :
                3
          :
             (X2[7:1] <= 44)?
              1
            :
              2
        :
           (X0[7:2] <= 29)?
             (X0[7:4] <= 7)?
              2
            :
              2
          :
            5
      :
        29
  :
     (X5[7:3] <= 3)?
       (X5[7:2] <= 8)?
         (X4[7:3] <= 23)?
          24
        :
           (X2[7:1] <= 43)?
            3
          :
            1
      :
        1
    :
      75
;
endmodule
