module tb();
