
`timescale 1ns/1ps
module top_tb();
`define EOF 32'hFFFF_FFFF
`define NULL 0
localparam period = 0;
localparam halfperiod = period/2;

reg [7:0] X0_reg;
reg [7:0] X1_reg;
reg [7:0] X4_reg;
reg [7:0] X9_reg;
reg [7:0] X12_reg;
reg [7:0] X28_reg;
reg [7:0] X30_reg;
reg [7:0] X32_reg;
reg [7:0] X37_reg;
reg [7:0] X38_reg;
reg [7:0] X41_reg;
reg [7:0] X42_reg;
reg [7:0] X44_reg;
reg [7:0] X49_reg;
reg [7:0] X51_reg;
reg [7:0] X52_reg;
reg [7:0] X54_reg;
reg [7:0] X55_reg;
reg [7:0] X56_reg;
reg [7:0] X57_reg;
reg [7:0] X58_reg;
reg [7:0] X62_reg;
reg [7:0] X63_reg;
reg [7:0] X65_reg;
reg [7:0] X69_reg;
reg [7:0] X73_reg;
reg [7:0] X90_reg;
reg [7:0] X93_reg;
reg [7:0] X101_reg;
reg [7:0] X102_reg;
reg [7:0] X106_reg;
reg [7:0] X113_reg;
reg [7:0] X114_reg;
reg [7:0] X115_reg;
reg [7:0] X118_reg;
reg [7:0] X125_reg;
reg [7:0] X128_reg;
reg [7:0] X133_reg;
reg [7:0] X136_reg;
reg [7:0] X137_reg;
reg [7:0] X139_reg;
reg [7:0] X141_reg;
reg [7:0] X142_reg;
reg [7:0] X147_reg;
reg [7:0] X148_reg;
reg [7:0] X155_reg;
reg [7:0] X159_reg;
reg [7:0] X161_reg;
reg [7:0] X162_reg;
reg [7:0] X165_reg;
reg [7:0] X169_reg;
reg [7:0] X170_reg;
reg [7:0] X172_reg;
reg [7:0] X180_reg;
reg [7:0] X181_reg;
reg [7:0] X185_reg;
reg [7:0] X190_reg;
reg [7:0] X192_reg;
reg [7:0] X198_reg;
reg [7:0] X199_reg;
reg [7:0] X209_reg;
reg [7:0] X210_reg;
reg [7:0] X227_reg;
reg [7:0] X238_reg;
reg [7:0] X240_reg;
reg [7:0] X244_reg;
reg [7:0] X245_reg;
reg [7:0] X248_reg;
reg [7:0] X258_reg;
reg [7:0] X259_reg;
reg [7:0] X263_reg;
reg [7:0] X265_reg;
reg [7:0] X268_reg;
reg [7:0] X270_reg;
reg [7:0] X273_reg;
reg [7:0] X274_reg;
reg [7:0] X275_reg;
reg [7:0] X276_reg;
reg [7:0] X283_reg;
reg [7:0] X286_reg;
reg [7:0] X287_reg;
reg [7:0] X290_reg;
reg [7:0] X296_reg;
reg [7:0] X300_reg;
reg [7:0] X301_reg;
reg [7:0] X302_reg;
reg [7:0] X310_reg;
reg [7:0] X312_reg;
reg [7:0] X313_reg;
reg [7:0] X319_reg;
reg [7:0] X320_reg;
reg [7:0] X323_reg;
reg [7:0] X324_reg;
reg [7:0] X326_reg;
reg [7:0] X327_reg;
reg [7:0] X330_reg;
reg [7:0] X331_reg;
reg [7:0] X335_reg;
reg [7:0] X336_reg;
reg [7:0] X340_reg;
reg [7:0] X342_reg;
reg [7:0] X358_reg;
reg [7:0] X361_reg;
reg [7:0] X362_reg;
reg [7:0] X370_reg;
reg [7:0] X371_reg;
reg [7:0] X376_reg;
reg [7:0] X380_reg;
reg [7:0] X387_reg;
reg [7:0] X388_reg;
reg [7:0] X394_reg;
reg [7:0] X395_reg;
reg [7:0] X403_reg;
reg [7:0] X405_reg;
reg [7:0] X409_reg;
reg [7:0] X410_reg;
reg [7:0] X414_reg;
reg [7:0] X428_reg;
reg [7:0] X432_reg;
reg [7:0] X434_reg;
reg [7:0] X435_reg;
reg [7:0] X445_reg;
reg [7:0] X449_reg;
reg [7:0] X452_reg;
reg [7:0] X455_reg;
reg [7:0] X457_reg;
reg [7:0] X458_reg;
reg [7:0] X460_reg;
reg [7:0] X462_reg;
reg [7:0] X477_reg;
reg [7:0] X481_reg;
reg [7:0] X483_reg;
reg [7:0] X488_reg;
reg [7:0] X489_reg;
reg [7:0] X498_reg;
reg [7:0] X504_reg;
reg [7:0] X509_reg;
reg [7:0] X514_reg;
reg [7:0] X524_reg;
reg [7:0] X527_reg;
reg [7:0] X535_reg;
reg [7:0] X537_reg;
reg [7:0] X539_reg;
reg [7:0] X542_reg;
reg [7:0] X550_reg;
reg [7:0] X554_reg;
reg [7:0] X558_reg;
reg [7:0] X560_reg;
wire [7:0] X0;
wire [7:0] X1;
wire [7:0] X4;
wire [7:0] X9;
wire [7:0] X12;
wire [7:0] X28;
wire [7:0] X30;
wire [7:0] X32;
wire [7:0] X37;
wire [7:0] X38;
wire [7:0] X41;
wire [7:0] X42;
wire [7:0] X44;
wire [7:0] X49;
wire [7:0] X51;
wire [7:0] X52;
wire [7:0] X54;
wire [7:0] X55;
wire [7:0] X56;
wire [7:0] X57;
wire [7:0] X58;
wire [7:0] X62;
wire [7:0] X63;
wire [7:0] X65;
wire [7:0] X69;
wire [7:0] X73;
wire [7:0] X90;
wire [7:0] X93;
wire [7:0] X101;
wire [7:0] X102;
wire [7:0] X106;
wire [7:0] X113;
wire [7:0] X114;
wire [7:0] X115;
wire [7:0] X118;
wire [7:0] X125;
wire [7:0] X128;
wire [7:0] X133;
wire [7:0] X136;
wire [7:0] X137;
wire [7:0] X139;
wire [7:0] X141;
wire [7:0] X142;
wire [7:0] X147;
wire [7:0] X148;
wire [7:0] X155;
wire [7:0] X159;
wire [7:0] X161;
wire [7:0] X162;
wire [7:0] X165;
wire [7:0] X169;
wire [7:0] X170;
wire [7:0] X172;
wire [7:0] X180;
wire [7:0] X181;
wire [7:0] X185;
wire [7:0] X190;
wire [7:0] X192;
wire [7:0] X198;
wire [7:0] X199;
wire [7:0] X209;
wire [7:0] X210;
wire [7:0] X227;
wire [7:0] X238;
wire [7:0] X240;
wire [7:0] X244;
wire [7:0] X245;
wire [7:0] X248;
wire [7:0] X258;
wire [7:0] X259;
wire [7:0] X263;
wire [7:0] X265;
wire [7:0] X268;
wire [7:0] X270;
wire [7:0] X273;
wire [7:0] X274;
wire [7:0] X275;
wire [7:0] X276;
wire [7:0] X283;
wire [7:0] X286;
wire [7:0] X287;
wire [7:0] X290;
wire [7:0] X296;
wire [7:0] X300;
wire [7:0] X301;
wire [7:0] X302;
wire [7:0] X310;
wire [7:0] X312;
wire [7:0] X313;
wire [7:0] X319;
wire [7:0] X320;
wire [7:0] X323;
wire [7:0] X324;
wire [7:0] X326;
wire [7:0] X327;
wire [7:0] X330;
wire [7:0] X331;
wire [7:0] X335;
wire [7:0] X336;
wire [7:0] X340;
wire [7:0] X342;
wire [7:0] X358;
wire [7:0] X361;
wire [7:0] X362;
wire [7:0] X370;
wire [7:0] X371;
wire [7:0] X376;
wire [7:0] X380;
wire [7:0] X387;
wire [7:0] X388;
wire [7:0] X394;
wire [7:0] X395;
wire [7:0] X403;
wire [7:0] X405;
wire [7:0] X409;
wire [7:0] X410;
wire [7:0] X414;
wire [7:0] X428;
wire [7:0] X432;
wire [7:0] X434;
wire [7:0] X435;
wire [7:0] X445;
wire [7:0] X449;
wire [7:0] X452;
wire [7:0] X455;
wire [7:0] X457;
wire [7:0] X458;
wire [7:0] X460;
wire [7:0] X462;
wire [7:0] X477;
wire [7:0] X481;
wire [7:0] X483;
wire [7:0] X488;
wire [7:0] X489;
wire [7:0] X498;
wire [7:0] X504;
wire [7:0] X509;
wire [7:0] X514;
wire [7:0] X524;
wire [7:0] X527;
wire [7:0] X535;
wire [7:0] X537;
wire [7:0] X539;
wire [7:0] X542;
wire [7:0] X550;
wire [7:0] X554;
wire [7:0] X558;
wire [7:0] X560;
wire [2:0] out;

integer fin, fout, r;

top DUT (X0, X1, X4, X9, X12, X28, X30, X32, X37, X38, X41, X42, X44, X49, X51, X52, X54, X55, X56, X57, X58, X62, X63, X65, X69, X73, X90, X93, X101, X102, X106, X113, X114, X115, X118, X125, X128, X133, X136, X137, X139, X141, X142, X147, X148, X155, X159, X161, X162, X165, X169, X170, X172, X180, X181, X185, X190, X192, X198, X199, X209, X210, X227, X238, X240, X244, X245, X248, X258, X259, X263, X265, X268, X270, X273, X274, X275, X276, X283, X286, X287, X290, X296, X300, X301, X302, X310, X312, X313, X319, X320, X323, X324, X326, X327, X330, X331, X335, X336, X340, X342, X358, X361, X362, X370, X371, X376, X380, X387, X388, X394, X395, X403, X405, X409, X410, X414, X428, X432, X434, X435, X445, X449, X452, X455, X457, X458, X460, X462, X477, X481, X483, X488, X489, X498, X504, X509, X514, X524, X527, X535, X537, X539, X542, X550, X554, X558, X560, out);

//read inp
initial begin
    $display($time, " << Starting the Simulation >>");
    fin = $fopen("/home/balkon00/PrintedTrees/test/pareto/sim/inputs.txt", "r");
    if (fin == `NULL) begin
        $display($time, " file not found");
        $finish;
    end
    fout = $fopen("/home/balkon00/PrintedTrees/test/pareto/sim/output.txt", "w");
    forever begin
        r = $fscanf(fin,"%d\t%d\t%d\t%d\t%d\t%d\t%d\t%d\t%d\t%d\t%d\t%d\t%d\t%d\t%d\t%d\t%d\t%d\t%d\t%d\t%d\t%d\t%d\t%d\t%d\t%d\t%d\t%d\t%d\t%d\t%d\t%d\t%d\t%d\t%d\t%d\t%d\t%d\t%d\t%d\t%d\t%d\t%d\t%d\t%d\t%d\t%d\t%d\t%d\t%d\t%d\t%d\t%d\t%d\t%d\t%d\t%d\t%d\t%d\t%d\t%d\t%d\t%d\t%d\t%d\t%d\t%d\t%d\t%d\t%d\t%d\t%d\t%d\t%d\t%d\t%d\t%d\t%d\t%d\t%d\t%d\t%d\t%d\t%d\t%d\t%d\t%d\t%d\t%d\t%d\t%d\t%d\t%d\t%d\t%d\t%d\t%d\t%d\t%d\t%d\t%d\t%d\t%d\t%d\t%d\t%d\t%d\t%d\t%d\t%d\t%d\t%d\t%d\t%d\t%d\t%d\t%d\t%d\t%d\t%d\t%d\t%d\t%d\t%d\t%d\t%d\t%d\t%d\t%d\t%d\t%d\t%d\t%d\t%d\t%d\t%d\t%d\t%d\t%d\t%d\t%d\t%d\t%d\t%d\t%d\t%d\t%d\t%d\n", X0_reg, X1_reg, X4_reg, X9_reg, X12_reg, X28_reg, X30_reg, X32_reg, X37_reg, X38_reg, X41_reg, X42_reg, X44_reg, X49_reg, X51_reg, X52_reg, X54_reg, X55_reg, X56_reg, X57_reg, X58_reg, X62_reg, X63_reg, X65_reg, X69_reg, X73_reg, X90_reg, X93_reg, X101_reg, X102_reg, X106_reg, X113_reg, X114_reg, X115_reg, X118_reg, X125_reg, X128_reg, X133_reg, X136_reg, X137_reg, X139_reg, X141_reg, X142_reg, X147_reg, X148_reg, X155_reg, X159_reg, X161_reg, X162_reg, X165_reg, X169_reg, X170_reg, X172_reg, X180_reg, X181_reg, X185_reg, X190_reg, X192_reg, X198_reg, X199_reg, X209_reg, X210_reg, X227_reg, X238_reg, X240_reg, X244_reg, X245_reg, X248_reg, X258_reg, X259_reg, X263_reg, X265_reg, X268_reg, X270_reg, X273_reg, X274_reg, X275_reg, X276_reg, X283_reg, X286_reg, X287_reg, X290_reg, X296_reg, X300_reg, X301_reg, X302_reg, X310_reg, X312_reg, X313_reg, X319_reg, X320_reg, X323_reg, X324_reg, X326_reg, X327_reg, X330_reg, X331_reg, X335_reg, X336_reg, X340_reg, X342_reg, X358_reg, X361_reg, X362_reg, X370_reg, X371_reg, X376_reg, X380_reg, X387_reg, X388_reg, X394_reg, X395_reg, X403_reg, X405_reg, X409_reg, X410_reg, X414_reg, X428_reg, X432_reg, X434_reg, X435_reg, X445_reg, X449_reg, X452_reg, X455_reg, X457_reg, X458_reg, X460_reg, X462_reg, X477_reg, X481_reg, X483_reg, X488_reg, X489_reg, X498_reg, X504_reg, X509_reg, X514_reg, X524_reg, X527_reg, X535_reg, X537_reg, X539_reg, X542_reg, X550_reg, X554_reg, X558_reg, X560_reg);
        #period $fwrite(fout, "%d\n", out);
        if ($feof(fin)) begin
            $display($time, " << Finishing the Simulation >>");
            $fclose(fin);
            $fclose(fout);
            $finish;
        end
    end
end

assign X0 = X0_reg;
assign X1 = X1_reg;
assign X4 = X4_reg;
assign X9 = X9_reg;
assign X12 = X12_reg;
assign X28 = X28_reg;
assign X30 = X30_reg;
assign X32 = X32_reg;
assign X37 = X37_reg;
assign X38 = X38_reg;
assign X41 = X41_reg;
assign X42 = X42_reg;
assign X44 = X44_reg;
assign X49 = X49_reg;
assign X51 = X51_reg;
assign X52 = X52_reg;
assign X54 = X54_reg;
assign X55 = X55_reg;
assign X56 = X56_reg;
assign X57 = X57_reg;
assign X58 = X58_reg;
assign X62 = X62_reg;
assign X63 = X63_reg;
assign X65 = X65_reg;
assign X69 = X69_reg;
assign X73 = X73_reg;
assign X90 = X90_reg;
assign X93 = X93_reg;
assign X101 = X101_reg;
assign X102 = X102_reg;
assign X106 = X106_reg;
assign X113 = X113_reg;
assign X114 = X114_reg;
assign X115 = X115_reg;
assign X118 = X118_reg;
assign X125 = X125_reg;
assign X128 = X128_reg;
assign X133 = X133_reg;
assign X136 = X136_reg;
assign X137 = X137_reg;
assign X139 = X139_reg;
assign X141 = X141_reg;
assign X142 = X142_reg;
assign X147 = X147_reg;
assign X148 = X148_reg;
assign X155 = X155_reg;
assign X159 = X159_reg;
assign X161 = X161_reg;
assign X162 = X162_reg;
assign X165 = X165_reg;
assign X169 = X169_reg;
assign X170 = X170_reg;
assign X172 = X172_reg;
assign X180 = X180_reg;
assign X181 = X181_reg;
assign X185 = X185_reg;
assign X190 = X190_reg;
assign X192 = X192_reg;
assign X198 = X198_reg;
assign X199 = X199_reg;
assign X209 = X209_reg;
assign X210 = X210_reg;
assign X227 = X227_reg;
assign X238 = X238_reg;
assign X240 = X240_reg;
assign X244 = X244_reg;
assign X245 = X245_reg;
assign X248 = X248_reg;
assign X258 = X258_reg;
assign X259 = X259_reg;
assign X263 = X263_reg;
assign X265 = X265_reg;
assign X268 = X268_reg;
assign X270 = X270_reg;
assign X273 = X273_reg;
assign X274 = X274_reg;
assign X275 = X275_reg;
assign X276 = X276_reg;
assign X283 = X283_reg;
assign X286 = X286_reg;
assign X287 = X287_reg;
assign X290 = X290_reg;
assign X296 = X296_reg;
assign X300 = X300_reg;
assign X301 = X301_reg;
assign X302 = X302_reg;
assign X310 = X310_reg;
assign X312 = X312_reg;
assign X313 = X313_reg;
assign X319 = X319_reg;
assign X320 = X320_reg;
assign X323 = X323_reg;
assign X324 = X324_reg;
assign X326 = X326_reg;
assign X327 = X327_reg;
assign X330 = X330_reg;
assign X331 = X331_reg;
assign X335 = X335_reg;
assign X336 = X336_reg;
assign X340 = X340_reg;
assign X342 = X342_reg;
assign X358 = X358_reg;
assign X361 = X361_reg;
assign X362 = X362_reg;
assign X370 = X370_reg;
assign X371 = X371_reg;
assign X376 = X376_reg;
assign X380 = X380_reg;
assign X387 = X387_reg;
assign X388 = X388_reg;
assign X394 = X394_reg;
assign X395 = X395_reg;
assign X403 = X403_reg;
assign X405 = X405_reg;
assign X409 = X409_reg;
assign X410 = X410_reg;
assign X414 = X414_reg;
assign X428 = X428_reg;
assign X432 = X432_reg;
assign X434 = X434_reg;
assign X435 = X435_reg;
assign X445 = X445_reg;
assign X449 = X449_reg;
assign X452 = X452_reg;
assign X455 = X455_reg;
assign X457 = X457_reg;
assign X458 = X458_reg;
assign X460 = X460_reg;
assign X462 = X462_reg;
assign X477 = X477_reg;
assign X481 = X481_reg;
assign X483 = X483_reg;
assign X488 = X488_reg;
assign X489 = X489_reg;
assign X498 = X498_reg;
assign X504 = X504_reg;
assign X509 = X509_reg;
assign X514 = X514_reg;
assign X524 = X524_reg;
assign X527 = X527_reg;
assign X535 = X535_reg;
assign X537 = X537_reg;
assign X539 = X539_reg;
assign X542 = X542_reg;
assign X550 = X550_reg;
assign X554 = X554_reg;
assign X558 = X558_reg;
assign X560 = X560_reg;

endmodule

