
`timescale 1ns/1ps
module top_tb();
`define EOF 32'hFFFF_FFFF
`define NULL 0
localparam period = 0;
localparam halfperiod = period/2;

reg [7:0] X2_reg;
reg [7:0] X6_reg;
reg [7:0] X9_reg;
reg [7:0] X10_reg;
reg [7:0] X12_reg;
reg [7:0] X14_reg;
reg [7:0] X23_reg;
reg [7:0] X28_reg;
reg [7:0] X32_reg;
reg [7:0] X36_reg;
reg [7:0] X37_reg;
reg [7:0] X40_reg;
reg [7:0] X41_reg;
reg [7:0] X42_reg;
reg [7:0] X43_reg;
reg [7:0] X50_reg;
reg [7:0] X51_reg;
reg [7:0] X54_reg;
reg [7:0] X55_reg;
reg [7:0] X56_reg;
reg [7:0] X57_reg;
reg [7:0] X58_reg;
reg [7:0] X63_reg;
reg [7:0] X65_reg;
reg [7:0] X68_reg;
reg [7:0] X69_reg;
reg [7:0] X74_reg;
reg [7:0] X76_reg;
reg [7:0] X77_reg;
reg [7:0] X86_reg;
reg [7:0] X88_reg;
reg [7:0] X89_reg;
reg [7:0] X100_reg;
reg [7:0] X102_reg;
reg [7:0] X111_reg;
reg [7:0] X115_reg;
reg [7:0] X117_reg;
reg [7:0] X118_reg;
reg [7:0] X128_reg;
reg [7:0] X131_reg;
reg [7:0] X133_reg;
reg [7:0] X139_reg;
reg [7:0] X140_reg;
reg [7:0] X141_reg;
reg [7:0] X144_reg;
reg [7:0] X145_reg;
reg [7:0] X147_reg;
reg [7:0] X150_reg;
reg [7:0] X152_reg;
reg [7:0] X158_reg;
reg [7:0] X175_reg;
reg [7:0] X178_reg;
reg [7:0] X179_reg;
reg [7:0] X181_reg;
reg [7:0] X185_reg;
reg [7:0] X187_reg;
reg [7:0] X189_reg;
reg [7:0] X196_reg;
reg [7:0] X197_reg;
reg [7:0] X198_reg;
reg [7:0] X203_reg;
reg [7:0] X204_reg;
reg [7:0] X214_reg;
reg [7:0] X221_reg;
reg [7:0] X224_reg;
reg [7:0] X230_reg;
reg [7:0] X238_reg;
reg [7:0] X243_reg;
reg [7:0] X246_reg;
reg [7:0] X252_reg;
reg [7:0] X257_reg;
reg [7:0] X264_reg;
reg [7:0] X266_reg;
reg [7:0] X270_reg;
reg [7:0] X276_reg;
reg [7:0] X280_reg;
reg [7:0] X288_reg;
reg [7:0] X293_reg;
reg [7:0] X295_reg;
reg [7:0] X300_reg;
reg [7:0] X301_reg;
reg [7:0] X302_reg;
reg [7:0] X305_reg;
reg [7:0] X306_reg;
reg [7:0] X317_reg;
reg [7:0] X321_reg;
reg [7:0] X330_reg;
reg [7:0] X331_reg;
reg [7:0] X335_reg;
reg [7:0] X339_reg;
reg [7:0] X343_reg;
reg [7:0] X357_reg;
reg [7:0] X358_reg;
reg [7:0] X365_reg;
reg [7:0] X369_reg;
reg [7:0] X371_reg;
reg [7:0] X374_reg;
reg [7:0] X387_reg;
reg [7:0] X390_reg;
reg [7:0] X394_reg;
reg [7:0] X396_reg;
reg [7:0] X407_reg;
reg [7:0] X410_reg;
reg [7:0] X415_reg;
reg [7:0] X417_reg;
reg [7:0] X418_reg;
reg [7:0] X427_reg;
reg [7:0] X434_reg;
reg [7:0] X435_reg;
reg [7:0] X440_reg;
reg [7:0] X448_reg;
reg [7:0] X449_reg;
reg [7:0] X453_reg;
reg [7:0] X454_reg;
reg [7:0] X464_reg;
reg [7:0] X467_reg;
reg [7:0] X476_reg;
reg [7:0] X485_reg;
reg [7:0] X486_reg;
reg [7:0] X490_reg;
reg [7:0] X491_reg;
reg [7:0] X492_reg;
reg [7:0] X494_reg;
reg [7:0] X498_reg;
reg [7:0] X504_reg;
reg [7:0] X507_reg;
reg [7:0] X509_reg;
reg [7:0] X510_reg;
reg [7:0] X515_reg;
reg [7:0] X536_reg;
reg [7:0] X546_reg;
reg [7:0] X552_reg;
reg [7:0] X554_reg;
reg [7:0] X555_reg;
reg [7:0] X557_reg;
reg [7:0] X558_reg;
reg [7:0] X559_reg;
reg [7:0] X560_reg;
wire [7:0] X2;
wire [7:0] X6;
wire [7:0] X9;
wire [7:0] X10;
wire [7:0] X12;
wire [7:0] X14;
wire [7:0] X23;
wire [7:0] X28;
wire [7:0] X32;
wire [7:0] X36;
wire [7:0] X37;
wire [7:0] X40;
wire [7:0] X41;
wire [7:0] X42;
wire [7:0] X43;
wire [7:0] X50;
wire [7:0] X51;
wire [7:0] X54;
wire [7:0] X55;
wire [7:0] X56;
wire [7:0] X57;
wire [7:0] X58;
wire [7:0] X63;
wire [7:0] X65;
wire [7:0] X68;
wire [7:0] X69;
wire [7:0] X74;
wire [7:0] X76;
wire [7:0] X77;
wire [7:0] X86;
wire [7:0] X88;
wire [7:0] X89;
wire [7:0] X100;
wire [7:0] X102;
wire [7:0] X111;
wire [7:0] X115;
wire [7:0] X117;
wire [7:0] X118;
wire [7:0] X128;
wire [7:0] X131;
wire [7:0] X133;
wire [7:0] X139;
wire [7:0] X140;
wire [7:0] X141;
wire [7:0] X144;
wire [7:0] X145;
wire [7:0] X147;
wire [7:0] X150;
wire [7:0] X152;
wire [7:0] X158;
wire [7:0] X175;
wire [7:0] X178;
wire [7:0] X179;
wire [7:0] X181;
wire [7:0] X185;
wire [7:0] X187;
wire [7:0] X189;
wire [7:0] X196;
wire [7:0] X197;
wire [7:0] X198;
wire [7:0] X203;
wire [7:0] X204;
wire [7:0] X214;
wire [7:0] X221;
wire [7:0] X224;
wire [7:0] X230;
wire [7:0] X238;
wire [7:0] X243;
wire [7:0] X246;
wire [7:0] X252;
wire [7:0] X257;
wire [7:0] X264;
wire [7:0] X266;
wire [7:0] X270;
wire [7:0] X276;
wire [7:0] X280;
wire [7:0] X288;
wire [7:0] X293;
wire [7:0] X295;
wire [7:0] X300;
wire [7:0] X301;
wire [7:0] X302;
wire [7:0] X305;
wire [7:0] X306;
wire [7:0] X317;
wire [7:0] X321;
wire [7:0] X330;
wire [7:0] X331;
wire [7:0] X335;
wire [7:0] X339;
wire [7:0] X343;
wire [7:0] X357;
wire [7:0] X358;
wire [7:0] X365;
wire [7:0] X369;
wire [7:0] X371;
wire [7:0] X374;
wire [7:0] X387;
wire [7:0] X390;
wire [7:0] X394;
wire [7:0] X396;
wire [7:0] X407;
wire [7:0] X410;
wire [7:0] X415;
wire [7:0] X417;
wire [7:0] X418;
wire [7:0] X427;
wire [7:0] X434;
wire [7:0] X435;
wire [7:0] X440;
wire [7:0] X448;
wire [7:0] X449;
wire [7:0] X453;
wire [7:0] X454;
wire [7:0] X464;
wire [7:0] X467;
wire [7:0] X476;
wire [7:0] X485;
wire [7:0] X486;
wire [7:0] X490;
wire [7:0] X491;
wire [7:0] X492;
wire [7:0] X494;
wire [7:0] X498;
wire [7:0] X504;
wire [7:0] X507;
wire [7:0] X509;
wire [7:0] X510;
wire [7:0] X515;
wire [7:0] X536;
wire [7:0] X546;
wire [7:0] X552;
wire [7:0] X554;
wire [7:0] X555;
wire [7:0] X557;
wire [7:0] X558;
wire [7:0] X559;
wire [7:0] X560;
wire [2:0] out;

integer fin, fout, r;

top DUT (X2, X6, X9, X10, X12, X14, X23, X28, X32, X36, X37, X40, X41, X42, X43, X50, X51, X54, X55, X56, X57, X58, X63, X65, X68, X69, X74, X76, X77, X86, X88, X89, X100, X102, X111, X115, X117, X118, X128, X131, X133, X139, X140, X141, X144, X145, X147, X150, X152, X158, X175, X178, X179, X181, X185, X187, X189, X196, X197, X198, X203, X204, X214, X221, X224, X230, X238, X243, X246, X252, X257, X264, X266, X270, X276, X280, X288, X293, X295, X300, X301, X302, X305, X306, X317, X321, X330, X331, X335, X339, X343, X357, X358, X365, X369, X371, X374, X387, X390, X394, X396, X407, X410, X415, X417, X418, X427, X434, X435, X440, X448, X449, X453, X454, X464, X467, X476, X485, X486, X490, X491, X492, X494, X498, X504, X507, X509, X510, X515, X536, X546, X552, X554, X555, X557, X558, X559, X560, out);

//read inp
initial begin
    $display($time, " << Starting the Simulation >>");
    fin = $fopen("/home/balkon00/PrintedTrees/test/pareto/sim/inputs.txt", "r");
    if (fin == `NULL) begin
        $display($time, " file not found");
        $finish;
    end
    fout = $fopen("/home/balkon00/PrintedTrees/test/pareto/sim/output.txt", "w");
    forever begin
        r = $fscanf(fin,"%d\t%d\t%d\t%d\t%d\t%d\t%d\t%d\t%d\t%d\t%d\t%d\t%d\t%d\t%d\t%d\t%d\t%d\t%d\t%d\t%d\t%d\t%d\t%d\t%d\t%d\t%d\t%d\t%d\t%d\t%d\t%d\t%d\t%d\t%d\t%d\t%d\t%d\t%d\t%d\t%d\t%d\t%d\t%d\t%d\t%d\t%d\t%d\t%d\t%d\t%d\t%d\t%d\t%d\t%d\t%d\t%d\t%d\t%d\t%d\t%d\t%d\t%d\t%d\t%d\t%d\t%d\t%d\t%d\t%d\t%d\t%d\t%d\t%d\t%d\t%d\t%d\t%d\t%d\t%d\t%d\t%d\t%d\t%d\t%d\t%d\t%d\t%d\t%d\t%d\t%d\t%d\t%d\t%d\t%d\t%d\t%d\t%d\t%d\t%d\t%d\t%d\t%d\t%d\t%d\t%d\t%d\t%d\t%d\t%d\t%d\t%d\t%d\t%d\t%d\t%d\t%d\t%d\t%d\t%d\t%d\t%d\t%d\t%d\t%d\t%d\t%d\t%d\t%d\t%d\t%d\t%d\t%d\t%d\t%d\t%d\t%d\t%d\n", X2_reg, X6_reg, X9_reg, X10_reg, X12_reg, X14_reg, X23_reg, X28_reg, X32_reg, X36_reg, X37_reg, X40_reg, X41_reg, X42_reg, X43_reg, X50_reg, X51_reg, X54_reg, X55_reg, X56_reg, X57_reg, X58_reg, X63_reg, X65_reg, X68_reg, X69_reg, X74_reg, X76_reg, X77_reg, X86_reg, X88_reg, X89_reg, X100_reg, X102_reg, X111_reg, X115_reg, X117_reg, X118_reg, X128_reg, X131_reg, X133_reg, X139_reg, X140_reg, X141_reg, X144_reg, X145_reg, X147_reg, X150_reg, X152_reg, X158_reg, X175_reg, X178_reg, X179_reg, X181_reg, X185_reg, X187_reg, X189_reg, X196_reg, X197_reg, X198_reg, X203_reg, X204_reg, X214_reg, X221_reg, X224_reg, X230_reg, X238_reg, X243_reg, X246_reg, X252_reg, X257_reg, X264_reg, X266_reg, X270_reg, X276_reg, X280_reg, X288_reg, X293_reg, X295_reg, X300_reg, X301_reg, X302_reg, X305_reg, X306_reg, X317_reg, X321_reg, X330_reg, X331_reg, X335_reg, X339_reg, X343_reg, X357_reg, X358_reg, X365_reg, X369_reg, X371_reg, X374_reg, X387_reg, X390_reg, X394_reg, X396_reg, X407_reg, X410_reg, X415_reg, X417_reg, X418_reg, X427_reg, X434_reg, X435_reg, X440_reg, X448_reg, X449_reg, X453_reg, X454_reg, X464_reg, X467_reg, X476_reg, X485_reg, X486_reg, X490_reg, X491_reg, X492_reg, X494_reg, X498_reg, X504_reg, X507_reg, X509_reg, X510_reg, X515_reg, X536_reg, X546_reg, X552_reg, X554_reg, X555_reg, X557_reg, X558_reg, X559_reg, X560_reg);
        #period $fwrite(fout, "%d\n", out);
        if ($feof(fin)) begin
            $display($time, " << Finishing the Simulation >>");
            $fclose(fin);
            $fclose(fout);
            $finish;
        end
    end
end

assign X2 = X2_reg;
assign X6 = X6_reg;
assign X9 = X9_reg;
assign X10 = X10_reg;
assign X12 = X12_reg;
assign X14 = X14_reg;
assign X23 = X23_reg;
assign X28 = X28_reg;
assign X32 = X32_reg;
assign X36 = X36_reg;
assign X37 = X37_reg;
assign X40 = X40_reg;
assign X41 = X41_reg;
assign X42 = X42_reg;
assign X43 = X43_reg;
assign X50 = X50_reg;
assign X51 = X51_reg;
assign X54 = X54_reg;
assign X55 = X55_reg;
assign X56 = X56_reg;
assign X57 = X57_reg;
assign X58 = X58_reg;
assign X63 = X63_reg;
assign X65 = X65_reg;
assign X68 = X68_reg;
assign X69 = X69_reg;
assign X74 = X74_reg;
assign X76 = X76_reg;
assign X77 = X77_reg;
assign X86 = X86_reg;
assign X88 = X88_reg;
assign X89 = X89_reg;
assign X100 = X100_reg;
assign X102 = X102_reg;
assign X111 = X111_reg;
assign X115 = X115_reg;
assign X117 = X117_reg;
assign X118 = X118_reg;
assign X128 = X128_reg;
assign X131 = X131_reg;
assign X133 = X133_reg;
assign X139 = X139_reg;
assign X140 = X140_reg;
assign X141 = X141_reg;
assign X144 = X144_reg;
assign X145 = X145_reg;
assign X147 = X147_reg;
assign X150 = X150_reg;
assign X152 = X152_reg;
assign X158 = X158_reg;
assign X175 = X175_reg;
assign X178 = X178_reg;
assign X179 = X179_reg;
assign X181 = X181_reg;
assign X185 = X185_reg;
assign X187 = X187_reg;
assign X189 = X189_reg;
assign X196 = X196_reg;
assign X197 = X197_reg;
assign X198 = X198_reg;
assign X203 = X203_reg;
assign X204 = X204_reg;
assign X214 = X214_reg;
assign X221 = X221_reg;
assign X224 = X224_reg;
assign X230 = X230_reg;
assign X238 = X238_reg;
assign X243 = X243_reg;
assign X246 = X246_reg;
assign X252 = X252_reg;
assign X257 = X257_reg;
assign X264 = X264_reg;
assign X266 = X266_reg;
assign X270 = X270_reg;
assign X276 = X276_reg;
assign X280 = X280_reg;
assign X288 = X288_reg;
assign X293 = X293_reg;
assign X295 = X295_reg;
assign X300 = X300_reg;
assign X301 = X301_reg;
assign X302 = X302_reg;
assign X305 = X305_reg;
assign X306 = X306_reg;
assign X317 = X317_reg;
assign X321 = X321_reg;
assign X330 = X330_reg;
assign X331 = X331_reg;
assign X335 = X335_reg;
assign X339 = X339_reg;
assign X343 = X343_reg;
assign X357 = X357_reg;
assign X358 = X358_reg;
assign X365 = X365_reg;
assign X369 = X369_reg;
assign X371 = X371_reg;
assign X374 = X374_reg;
assign X387 = X387_reg;
assign X390 = X390_reg;
assign X394 = X394_reg;
assign X396 = X396_reg;
assign X407 = X407_reg;
assign X410 = X410_reg;
assign X415 = X415_reg;
assign X417 = X417_reg;
assign X418 = X418_reg;
assign X427 = X427_reg;
assign X434 = X434_reg;
assign X435 = X435_reg;
assign X440 = X440_reg;
assign X448 = X448_reg;
assign X449 = X449_reg;
assign X453 = X453_reg;
assign X454 = X454_reg;
assign X464 = X464_reg;
assign X467 = X467_reg;
assign X476 = X476_reg;
assign X485 = X485_reg;
assign X486 = X486_reg;
assign X490 = X490_reg;
assign X491 = X491_reg;
assign X492 = X492_reg;
assign X494 = X494_reg;
assign X498 = X498_reg;
assign X504 = X504_reg;
assign X507 = X507_reg;
assign X509 = X509_reg;
assign X510 = X510_reg;
assign X515 = X515_reg;
assign X536 = X536_reg;
assign X546 = X546_reg;
assign X552 = X552_reg;
assign X554 = X554_reg;
assign X555 = X555_reg;
assign X557 = X557_reg;
assign X558 = X558_reg;
assign X559 = X559_reg;
assign X560 = X560_reg;

endmodule

