module top(X0, X4, X12, X13, X39, X55, X74, X88, X91, X101, X110, X112, X124, X135, X161, X165, X170, X180, X195, X205, X206, X215, X218, X220, X221, X226, X229, X234, X235, X240, X246, X257, X264, X267, X275, X276, out);
input [7:0] X0;
input [7:0] X4;
input [7:0] X12;
input [7:0] X13;
input [7:0] X39;
input [7:0] X55;
input [7:0] X74;
input [7:0] X88;
input [7:0] X91;
input [7:0] X101;
input [7:0] X110;
input [7:0] X112;
input [7:0] X124;
input [7:0] X135;
input [7:0] X161;
input [7:0] X165;
input [7:0] X170;
input [7:0] X180;
input [7:0] X195;
input [7:0] X205;
input [7:0] X206;
input [7:0] X215;
input [7:0] X218;
input [7:0] X220;
input [7:0] X221;
input [7:0] X226;
input [7:0] X229;
input [7:0] X234;
input [7:0] X235;
input [7:0] X240;
input [7:0] X246;
input [7:0] X257;
input [7:0] X264;
input [7:0] X267;
input [7:0] X275;
input [7:0] X276;
output [4:0] out;
assign out = 
   (X195 <= 81)?
     (X13 <= 31)?
       (X226 <= 109)?
         (X264 <= 107)?
          14
        :
           (X275 <= 167)?
            3
          :
            2
      :
         (X161 <= 217)?
          3
        :
          1
    :
       (X226 <= 111)?
         (X110 <= 61)?
           (X205 <= 138)?
             (X234 <= 103)?
               (X135 <= 94)?
                3
              :
                3
            :
               (X246 <= 132)?
                 (X4 <= 131)?
                  1
                :
                  1
              :
                7
          :
             (X180 <= 153)?
               (X101 <= 64)?
                 (X124 <= 103)?
                  117
                :
                   (X91 <= 97)?
                     (X0 <= 222)?
                      21
                    :
                       (X55 <= 61)?
                        1
                      :
                        1
                  :
                    2
              :
                 (X215 <= 140)?
                  2
                :
                  3
            :
              2
        :
           (X267 <= 125)?
            4
          :
             (X229 <= 254)?
              1
            :
              1
      :
         (X13 <= 109)?
           (X88 <= 93)?
             (X39 <= 66)?
               (X161 <= 186)?
                1
              :
                2
            :
               (X218 <= 66)?
                10
              :
                1
          :
             (X170 <= 189)?
              6
            :
              1
        :
           (X12 <= 149)?
            1
          :
            6
  :
     (X240 <= 14)?
       (X220 <= 12)?
        8
      :
        2
    :
       (X112 <= 151)?
         (X74 <= 81)?
           (X275 <= 116)?
             (X13 <= 43)?
               (X206 <= 73)?
                1
              :
                2
            :
              14
          :
             (X13 <= 120)?
               (X257 <= 122)?
                 (X221 <= 196)?
                  3
                :
                  5
              :
                17
            :
               (X276 <= 123)?
                2
              :
                1
        :
           (X235 <= 118)?
             (X165 <= 178)?
              2
            :
              1
          :
            7
      :
         (X226 <= 90)?
          7
        :
          1
;
endmodule
