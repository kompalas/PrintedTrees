module top(X0, X1, X2, X3, X4, X5, X6, X7, X8, X9, X10, out);
input [7:0] X0;
input [7:0] X1;
input [7:0] X2;
input [7:0] X3;
input [7:0] X4;
input [7:0] X5;
input [7:0] X6;
input [7:0] X7;
input [7:0] X8;
input [7:0] X9;
input [7:0] X10;
output [3:0] out;
assign out = 
   (X10[7:3] <= 11)?
     (X0 <= 136)?
       (X6[7:2] <= 20)?
         (X9[7:1] <= 17)?
           (X3[7:5] <= 5)?
             (X4[7:2] <= 6)?
               (X6[7:3] <= 11)?
                 (X2 <= 84)?
                   (X9[7:2] <= 9)?
                     (X0[7:1] <= 42)?
                       (X9[7:4] <= 3)?
                        13
                      :
                         (X0[7:5] <= 2)?
                           (X4[7:1] <= 17)?
                            1
                          :
                            5
                        :
                          2
                    :
                       (X10[7:1] <= 29)?
                        1
                      :
                        2
                  :
                    20
                :
                   (X1[7:4] <= 4)?
                    1
                  :
                     (X9 <= 23)?
                      1
                    :
                      4
              :
                3
            :
               (X4[7:2] <= 20)?
                 (X7 <= 139)?
                  20
                :
                   (X7[7:2] <= 36)?
                     (X0[7:3] <= 11)?
                      2
                    :
                      3
                  :
                    12
              :
                1
          :
             (X2[7:1] <= 17)?
              1
            :
              3
        :
           (X1[7:1] <= 48)?
             (X1[7:2] <= 5)?
              5
            :
               (X0[7:3] <= 13)?
                 (X1 <= 47)?
                   (X7[7:2] <= 29)?
                    3
                  :
                     (X6[7:3] <= 12)?
                       (X1[7:3] <= 11)?
                        7
                      :
                         (X10[7:4] <= 5)?
                          1
                        :
                          1
                    :
                      1
                :
                   (X0[7:1] <= 24)?
                    11
                  :
                     (X2[7:4] <= 0)?
                      8
                    :
                       (X6[7:1] <= 16)?
                         (X7[7:4] <= 7)?
                          7
                        :
                           (X7[7:3] <= 20)?
                             (X0[7:4] <= 4)?
                               (X4[7:4] <= 4)?
                                 (X8[7:1] <= 57)?
                                  11
                                :
                                   (X8[7:2] <= 33)?
                                    3
                                  :
                                     (X10[7:3] <= 6)?
                                      1
                                    :
                                       (X9[7:2] <= 14)?
                                        1
                                      :
                                        7
                              :
                                2
                            :
                              3
                          :
                             (X8[7:3] <= 14)?
                               (X7[7:2] <= 36)?
                                1
                              :
                                1
                            :
                              8
                      :
                         (X3[7:5] <= 1)?
                          14
                        :
                           (X0[7:2] <= 18)?
                             (X4[7:2] <= 8)?
                               (X4[7:1] <= 17)?
                                 (X1[7:2] <= 14)?
                                  1
                                :
                                  13
                              :
                                 (X1 <= 83)?
                                   (X2[7:4] <= 9)?
                                     (X1[7:2] <= 17)?
                                      2
                                    :
                                       (X0[7:1] <= 37)?
                                        3
                                      :
                                        1
                                  :
                                    4
                                :
                                  7
                            :
                              10
                          :
                             (X9[7:4] <= 2)?
                              1
                            :
                              8
              :
                 (X0[7:1] <= 62)?
                   (X9[7:2] <= 14)?
                     (X9[7:3] <= 8)?
                      18
                    :
                       (X0[7:2] <= 31)?
                        1
                      :
                        1
                  :
                     (X0[7:2] <= 24)?
                       (X9 <= 51)?
                        3
                      :
                         (X9[7:2] <= 41)?
                          7
                        :
                          1
                    :
                       (X7[7:2] <= 55)?
                        13
                      :
                         (X1[7:1] <= 34)?
                          1
                        :
                          2
                :
                   (X2[7:1] <= 66)?
                     (X0 <= 133)?
                      7
                    :
                      1
                  :
                    5
          :
             (X10[7:1] <= 18)?
              2
            :
               (X1[7:3] <= 17)?
                 (X0 <= 101)?
                   (X8[7:2] <= 27)?
                     (X5[7:2] <= 11)?
                       (X10[7:5] <= 3)?
                        2
                      :
                        1
                    :
                      8
                  :
                     (X7[7:3] <= 16)?
                       (X9[7:2] <= 6)?
                         (X5[7:2] <= 8)?
                          2
                        :
                          3
                      :
                         (X0[7:1] <= 26)?
                           (X4[7:4] <= 4)?
                             (X7[7:4] <= 7)?
                              6
                            :
                              1
                          :
                            2
                        :
                          13
                    :
                      13
                :
                   (X10[7:1] <= 24)?
                    3
                  :
                     (X2[7:1] <= 16)?
                      1
                    :
                      1
              :
                 (X9[7:3] <= 9)?
                  2
                :
                  2
      :
         (X4[7:2] <= 5)?
           (X6[7:3] <= 15)?
            2
          :
            3
        :
          45
    :
       (X9[7:2] <= 12)?
         (X1[7:3] <= 10)?
          5
        :
          1
      :
         (X5[7:2] <= 16)?
           (X9[7:5] <= 4)?
            13
          :
             (X0[7:3] <= 25)?
               (X9[7:2] <= 21)?
                1
              :
                3
            :
               (X7[7:4] <= 12)?
                1
              :
                2
        :
          2
  :
     (X9[7:2] <= 15)?
       (X10[7:3] <= 16)?
         (X6[7:2] <= 6)?
           (X1[7:4] <= 7)?
             (X3[7:3] <= 2)?
               (X8[7:4] <= 11)?
                 (X7[7:2] <= 29)?
                  5
                :
                   (X8[7:2] <= 22)?
                    1
                  :
                    2
              :
                 (X2[7:2] <= 1)?
                   (X8[7:4] <= 8)?
                    2
                  :
                     (X3[7:3] <= 2)?
                      1
                    :
                      1
                :
                  7
            :
               (X9[7:1] <= 19)?
                 (X1[7:4] <= 5)?
                   (X3 <= 23)?
                    5
                  :
                     (X0[7:2] <= 17)?
                       (X9[7:3] <= 4)?
                        4
                      :
                        2
                    :
                       (X0[7:3] <= 9)?
                        4
                      :
                         (X8[7:2] <= 27)?
                          6
                        :
                          1
                :
                   (X4[7:4] <= 5)?
                     (X6[7:2] <= 2)?
                      1
                    :
                       (X5[7:5] <= 3)?
                        15
                      :
                        1
                  :
                    1
              :
                 (X4[7:2] <= 7)?
                   (X10[7:3] <= 13)?
                    4
                  :
                     (X0[7:2] <= 27)?
                      1
                    :
                      1
                :
                   (X0[7:2] <= 36)?
                     (X6[7:2] <= 5)?
                      9
                    :
                      1
                  :
                    1
          :
             (X9[7:1] <= 15)?
               (X6[7:4] <= 4)?
                 (X1[7:4] <= 13)?
                   (X1[7:4] <= 8)?
                    1
                  :
                    3
                :
                  2
              :
                1
            :
               (X2[7:4] <= 2)?
                3
              :
                 (X7[7:3] <= 19)?
                  3
                :
                  1
        :
           (X9[7:3] <= 5)?
             (X10[7:1] <= 54)?
               (X3[7:2] <= 11)?
                 (X3[7:3] <= 6)?
                   (X4[7:4] <= 4)?
                    4
                  :
                    8
                :
                  25
              :
                 (X10[7:3] <= 11)?
                  2
                :
                  4
            :
               (X5[7:2] <= 20)?
                 (X2[7:3] <= 3)?
                   (X2[7:2] <= 1)?
                    1
                  :
                    2
                :
                  2
              :
                1
          :
             (X7[7:1] <= 76)?
               (X0[7:2] <= 23)?
                 (X1[7:1] <= 26)?
                   (X10[7:1] <= 33)?
                    1
                  :
                    4
                :
                   (X2[7:2] <= 5)?
                     (X5 <= 123)?
                       (X0[7:2] <= 21)?
                        19
                      :
                        1
                    :
                      2
                  :
                     (X2[7:3] <= 12)?
                       (X9[7:2] <= 10)?
                        8
                      :
                         (X6[7:3] <= 6)?
                          1
                        :
                          2
                    :
                       (X9[7:1] <= 25)?
                         (X5[7:4] <= 4)?
                           (X3[7:1] <= 15)?
                            4
                          :
                            3
                        :
                          9
                      :
                        2
              :
                 (X0[7:3] <= 14)?
                  1
                :
                  6
            :
              10
      :
         (X1[7:2] <= 18)?
           (X3[7:3] <= 9)?
             (X2[7:2] <= 44)?
               (X0[7:2] <= 3)?
                1
              :
                 (X4[7:1] <= 4)?
                  2
                :
                   (X6[7:4] <= 1)?
                     (X0[7:4] <= 9)?
                       (X0[7:4] <= 5)?
                         (X6[7:2] <= 3)?
                          1
                        :
                           (X6[7:4] <= 2)?
                            9
                          :
                             (X7[7:3] <= 13)?
                              1
                            :
                              1
                      :
                        3
                    :
                      8
                  :
                    20
            :
               (X8[7:2] <= 25)?
                1
              :
                1
          :
             (X2[7:2] <= 27)?
               (X7[7:5] <= 3)?
                1
              :
                2
            :
              5
        :
           (X7[7:2] <= 18)?
             (X8[7:1] <= 108)?
               (X2[7:3] <= 1)?
                 (X9 <= 33)?
                  3
                :
                  2
              :
                6
            :
              2
          :
             (X1[7:2] <= 33)?
               (X1 <= 84)?
                1
              :
                 (X4[7:3] <= 2)?
                  1
                :
                  7
            :
               (X1[7:5] <= 5)?
                1
              :
                1
    :
       (X10[7:2] <= 32)?
         (X1[7:1] <= 24)?
           (X6[7:3] <= 9)?
             (X8[7:3] <= 16)?
               (X0[7:3] <= 10)?
                 (X7[7:3] <= 13)?
                   (X10[7:3] <= 18)?
                    1
                  :
                    1
                :
                  2
              :
                 (X2[7:1] <= 83)?
                   (X3[7:2] <= 12)?
                     (X3[7:2] <= 10)?
                       (X6[7:2] <= 4)?
                         (X10[7:2] <= 21)?
                          7
                        :
                           (X1[7:2] <= 9)?
                            1
                          :
                            3
                      :
                         (X0[7:1] <= 53)?
                          3
                        :
                           (X7 <= 163)?
                             (X7[7:4] <= 7)?
                               (X2[7:2] <= 30)?
                                3
                              :
                                2
                            :
                              11
                          :
                            1
                    :
                       (X8[7:3] <= 9)?
                        1
                      :
                        1
                  :
                    6
                :
                  5
            :
               (X5[7:3] <= 5)?
                 (X9[7:2] <= 19)?
                   (X2[7:2] <= 23)?
                    3
                  :
                     (X2[7:4] <= 9)?
                       (X6[7:3] <= 1)?
                        1
                      :
                         (X6[7:3] <= 2)?
                           (X4[7:3] <= 3)?
                            2
                          :
                            1
                        :
                          2
                    :
                      5
                :
                   (X2[7:2] <= 37)?
                    8
                  :
                    1
              :
                 (X9[7:4] <= 7)?
                  10
                :
                   (X7[7:2] <= 27)?
                    5
                  :
                     (X7[7:4] <= 10)?
                       (X1[7:4] <= 4)?
                         (X10[7:2] <= 22)?
                          2
                        :
                          2
                      :
                        6
                    :
                      2
          :
             (X5[7:2] <= 30)?
               (X2[7:2] <= 36)?
                 (X8[7:3] <= 15)?
                  8
                :
                   (X2[7:2] <= 29)?
                    5
                  :
                    2
              :
                3
            :
               (X0[7:2] <= 20)?
                4
              :
                5
        :
           (X6[7:1] <= 36)?
             (X4[7:4] <= 2)?
               (X1[7:2] <= 26)?
                 (X1[7:2] <= 16)?
                   (X7[7:1] <= 68)?
                     (X7[7:4] <= 9)?
                       (X9[7:2] <= 18)?
                        8
                      :
                         (X7[7:4] <= 6)?
                          2
                        :
                          1
                    :
                      2
                  :
                     (X9[7:2] <= 14)?
                      1
                    :
                      12
                :
                   (X0[7:4] <= 3)?
                     (X8[7:2] <= 48)?
                      17
                    :
                      1
                  :
                     (X1[7:1] <= 33)?
                      3
                    :
                       (X8[7:4] <= 4)?
                        3
                      :
                         (X8[7:5] <= 7)?
                          20
                        :
                           (X2[7:3] <= 0)?
                            6
                          :
                            6
              :
                 (X1[7:3] <= 11)?
                  4
                :
                   (X10[7:3] <= 14)?
                     (X7[7:3] <= 22)?
                      5
                    :
                      3
                  :
                     (X1[7:1] <= 68)?
                      11
                    :
                      1
            :
               (X6[7:2] <= 14)?
                 (X2[7:2] <= 14)?
                   (X3 <= 26)?
                    2
                  :
                     (X3[7:1] <= 27)?
                       (X3[7:2] <= 9)?
                        4
                      :
                         (X5[7:2] <= 23)?
                          1
                        :
                          1
                    :
                      1
                :
                   (X2[7:3] <= 20)?
                     (X4[7:4] <= 3)?
                      12
                    :
                      1
                  :
                    2
              :
                6
          :
             (X9[7:2] <= 34)?
               (X2[7:3] <= 7)?
                 (X3[7:1] <= 13)?
                  1
                :
                   (X10[7:1] <= 56)?
                    1
                  :
                    1
              :
                15
            :
              4
      :
         (X10[7:4] <= 13)?
           (X9[7:1] <= 28)?
             (X6 <= 9)?
               (X3[7:4] <= 4)?
                1
              :
                6
            :
               (X3[7:2] <= 7)?
                 (X2[7:3] <= 16)?
                  1
                :
                  1
              :
                 (X0[7:1] <= 90)?
                   (X9[7:5] <= 5)?
                    14
                  :
                    1
                :
                  1
          :
             (X5[7:4] <= 6)?
               (X9[7:4] <= 6)?
                 (X0[7:1] <= 62)?
                  22
                :
                   (X3[7:3] <= 4)?
                    1
                  :
                    3
              :
                 (X5[7:2] <= 6)?
                   (X1[7:2] <= 14)?
                    1
                  :
                    5
                :
                  3
            :
               (X3[7:2] <= 10)?
                 (X10[7:5] <= 8)?
                  4
                :
                   (X2 <= 16)?
                    3
                  :
                     (X6[7:1] <= 14)?
                      4
                    :
                       (X6[7:1] <= 17)?
                        3
                      :
                         (X4[7:2] <= 2)?
                          2
                        :
                           (X8[7:3] <= 15)?
                             (X10[7:3] <= 19)?
                              2
                            :
                               (X4[7:3] <= 8)?
                                2
                              :
                                1
                          :
                            6
              :
                 (X10[7:1] <= 87)?
                  3
                :
                  1
        :
           (X6[7:1] <= 21)?
             (X4[7:2] <= 6)?
              2
            :
               (X9 <= 67)?
                3
              :
                2
          :
             (X5[7:4] <= 4)?
              2
            :
              3
;
endmodule
