module top(X13, X27, X235, X264, X278, out);
input [7:0] X13;
input [7:0] X27;
input [7:0] X235;
input [7:0] X264;
input [7:0] X278;
output [4:0] out;
assign out = 
   (X278 <= 9)?
    167
  :
     (X278 <= 26)?
      24
    :
       (X278 <= 145)?
         (X13 <= 33)?
           (X27 <= 190)?
            17
          :
            1
        :
           (X278 <= 43)?
            11
          :
             (X278 <= 60)?
              7
            :
               (X278 <= 85)?
                9
              :
                 (X235 <= 146)?
                   (X264 <= 114)?
                    2
                  :
                    1
                :
                  6
      :
         (X278 <= 188)?
          33
        :
           (X278 <= 239)?
            4
          :
            12
;
endmodule
