module top(X0, X1, X2, X3, X4, X5, X6, X7, X8, X9, X10, X11, X12, X13, X14, X15, out);
input [7:0] X0;
input [7:0] X1;
input [7:0] X2;
input [7:0] X3;
input [7:0] X4;
input [7:0] X5;
input [7:0] X6;
input [7:0] X7;
input [7:0] X8;
input [7:0] X9;
input [7:0] X10;
input [7:0] X11;
input [7:0] X12;
input [7:0] X13;
input [7:0] X14;
input [7:0] X15;
output [3:0] out;
assign out = 
   (X15[7:5] <= 0)?
     (X4[7:6] <= 1)?
       (X9[7:6] <= 0)?
         (X14[7:6] <= 0)?
          349
        :
           (X13[7:6] <= 0)?
             (X12[7:3] <= 15)?
              19
            :
              21
          :
             (X9[7:6] <= 0)?
              1
            :
              28
      :
         (X5[7:5] <= 0)?
           (X7[7:5] <= 5)?
             (X15[7:6] <= 0)?
               (X5[7:5] <= 0)?
                2
              :
                 (X9[7:5] <= 5)?
                  682
                :
                   (X11[7:6] <= 0)?
                    1
                  :
                    8
            :
               (X5[7:5] <= 0)?
                17
              :
                2
          :
             (X10[7:4] <= 11)?
               (X0[7:5] <= 5)?
                 (X13[7:5] <= 0)?
                   (X12[7:6] <= 0)?
                    1
                  :
                    1
                :
                  21
              :
                 (X13[7:5] <= 0)?
                  4
                :
                  1
            :
              38
        :
           (X9[7:6] <= 2)?
             (X14[7:5] <= 0)?
               (X6[7:6] <= 0)?
                 (X10[7:6] <= 0)?
                   (X7[7:6] <= 0)?
                    1
                  :
                    4
                :
                   (X2[7:6] <= 0)?
                     (X0[7:5] <= 0)?
                      2
                    :
                       (X5[7:6] <= 0)?
                        1
                      :
                        1
                  :
                     (X1[7:6] <= 1)?
                      1
                    :
                      91
              :
                 (X9[7:6] <= 0)?
                   (X0[7:5] <= 5)?
                    1
                  :
                    7
                :
                  33
            :
               (X10[7:6] <= 2)?
                 (X12[7:6] <= 3)?
                  19
                :
                   (X7[7:5] <= 3)?
                    6
                  :
                    1
              :
                 (X9[7:5] <= 2)?
                   (X13[7:6] <= 0)?
                     (X8[7:6] <= 0)?
                       (X6[7:6] <= 0)?
                        1
                      :
                        1
                    :
                      3
                  :
                    56
                :
                   (X5[7:4] <= 8)?
                    2
                  :
                    7
          :
             (X0[7:6] <= 0)?
               (X7[7:6] <= 4)?
                 (X11[7:6] <= 0)?
                   (X3[7:6] <= 3)?
                    1
                  :
                    3
                :
                  3
              :
                 (X1[7:5] <= 0)?
                  3
                :
                  24
            :
               (X1[7:6] <= 2)?
                207
              :
                 (X7[7:5] <= 1)?
                   (X13[7:5] <= 1)?
                    1
                  :
                    5
                :
                   (X5[7:6] <= 4)?
                    29
                  :
                    2
    :
       (X14[7:6] <= 0)?
         (X3[7:6] <= 4)?
           (X10[7:5] <= 4)?
             (X7[7:6] <= 2)?
               (X9[7:4] <= 4)?
                13
              :
                 (X5[7:6] <= 0)?
                  11
                :
                  1
            :
               (X0[7:6] <= 0)?
                 (X8[7:6] <= 0)?
                   (X13[7:5] <= 0)?
                     (X12[7:6] <= 0)?
                      1
                    :
                       (X1[7:6] <= 0)?
                        1
                      :
                        1
                  :
                    6
                :
                   (X3[7:5] <= 3)?
                     (X2[7:6] <= 0)?
                       (X3[7:6] <= 1)?
                         (X4[7:6] <= 0)?
                          5
                        :
                          1
                      :
                        2
                    :
                       (X13[7:4] <= 4)?
                        211
                      :
                        1
                  :
                     (X2[7:6] <= 0)?
                      9
                    :
                      4
              :
                 (X10[7:6] <= 0)?
                   (X3[7:5] <= 2)?
                     (X5[7:6] <= 1)?
                      2
                    :
                       (X5[7:6] <= 2)?
                        1
                      :
                        1
                  :
                    43
                :
                   (X0[7:5] <= 0)?
                     (X9[7:6] <= 0)?
                      5
                    :
                       (X3[7:6] <= 2)?
                         (X2[7:5] <= 0)?
                          1
                        :
                          1
                      :
                        3
                  :
                     (X7[7:6] <= 1)?
                      1
                    :
                      29
          :
             (X1[7:5] <= 0)?
               (X6[7:6] <= 0)?
                 (X13[7:5] <= 0)?
                  6
                :
                  4
              :
                11
            :
               (X9[7:6] <= 0)?
                 (X0[7:5] <= 1)?
                  2
                :
                  3
              :
                 (X0[7:5] <= 0)?
                   (X3[7:6] <= 0)?
                    10
                  :
                     (X2[7:6] <= 0)?
                      3
                    :
                       (X2[7:5] <= 3)?
                        2
                      :
                        1
                :
                   (X9[7:6] <= 0)?
                     (X0[7:6] <= 0)?
                      2
                    :
                      5
                  :
                    163
        :
           (X7[7:6] <= 3)?
             (X2[7:5] <= 5)?
               (X4[7:6] <= 0)?
                 (X9[7:6] <= 0)?
                   (X0[7:6] <= 1)?
                    2
                  :
                    7
                :
                   (X6[7:5] <= 4)?
                     (X2[7:5] <= 0)?
                      6
                    :
                       (X14[7:6] <= 1)?
                         (X1[7:6] <= 0)?
                          1
                        :
                           (X10[7:6] <= 0)?
                            1
                          :
                            23
                      :
                        2
                  :
                    9
              :
                 (X12[7:6] <= 0)?
                   (X15[7:5] <= 0)?
                    6
                  :
                     (X13[7:6] <= 0)?
                      1
                    :
                      3
                :
                   (X9[7:5] <= 0)?
                     (X15[7:6] <= 0)?
                      3
                    :
                       (X14[7:6] <= 0)?
                        1
                      :
                        2
                  :
                     (X3[7:4] <= 13)?
                       (X0[7:6] <= 0)?
                         (X6[7:6] <= 1)?
                           (X6[7:6] <= 1)?
                            1
                          :
                            16
                        :
                           (X1[7:5] <= 3)?
                            2
                          :
                            3
                      :
                         (X1[7:6] <= 0)?
                          1
                        :
                          3
                    :
                       (X5[7:4] <= 7)?
                        1
                      :
                         (X13[7:5] <= 0)?
                           (X2[7:6] <= 1)?
                            643
                          :
                             (X13[7:6] <= 0)?
                              16
                            :
                              1
                        :
                           (X10[7:6] <= 0)?
                            1
                          :
                            1
            :
               (X5[7:6] <= 2)?
                 (X13[7:5] <= 0)?
                   (X4[7:5] <= 2)?
                     (X2[7:5] <= 5)?
                      2
                    :
                      9
                  :
                     (X10[7:6] <= 0)?
                      2
                    :
                      23
                :
                   (X9[7:5] <= 0)?
                     (X9[7:6] <= 1)?
                      11
                    :
                      1
                  :
                    20
              :
                 (X1[7:6] <= 0)?
                  8
                :
                   (X6[7:5] <= 2)?
                     (X11[7:6] <= 0)?
                      64
                    :
                      1
                  :
                     (X15[7:6] <= 0)?
                       (X11[7:5] <= 1)?
                        1
                      :
                        2
                    :
                      2
          :
             (X5[7:6] <= 2)?
              92
            :
               (X2[7:6] <= 0)?
                 (X11[7:6] <= 0)?
                   (X10[7:6] <= 0)?
                    2
                  :
                    25
                :
                   (X2[7:6] <= 0)?
                    55
                  :
                     (X1[7:6] <= 3)?
                       (X1[7:6] <= 0)?
                        1
                      :
                         (X14[7:6] <= 1)?
                          1
                        :
                          1
                    :
                      4
              :
                 (X13[7:6] <= 0)?
                   (X11[7:6] <= 0)?
                    1
                  :
                    76
                :
                   (X11[7:5] <= 1)?
                    2
                  :
                    1
      :
         (X3[7:5] <= 3)?
           (X6[7:5] <= 0)?
             (X9[7:5] <= 0)?
               (X14[7:5] <= 6)?
                1
              :
                1
            :
              38
          :
             (X8[7:5] <= 0)?
               (X8[7:6] <= 2)?
                6
              :
                1
            :
               (X1[7:6] <= 1)?
                 (X10[7:4] <= 0)?
                   (X6[7:6] <= 0)?
                    12
                  :
                    4
                :
                   (X13[7:5] <= 0)?
                    257
                  :
                    1
              :
                 (X14[7:4] <= 13)?
                  3
                :
                  1
        :
           (X8[7:6] <= 0)?
             (X9[7:6] <= 0)?
               (X8[7:6] <= 0)?
                 (X4[7:6] <= 0)?
                   (X0[7:6] <= 0)?
                    15
                  :
                     (X5[7:6] <= 2)?
                      4
                    :
                      4
                :
                  105
              :
                 (X4[7:6] <= 0)?
                   (X8[7:5] <= 1)?
                     (X7[7:6] <= 0)?
                       (X12[7:6] <= 0)?
                        1
                      :
                        2
                    :
                       (X7[7:6] <= 1)?
                        7
                      :
                        1
                  :
                    15
                :
                   (X1[7:5] <= 3)?
                    26
                  :
                     (X6[7:5] <= 1)?
                      3
                    :
                      1
            :
               (X9[7:4] <= 7)?
                 (X5[7:4] <= 11)?
                  335
                :
                   (X2[7:6] <= 0)?
                    56
                  :
                     (X4[7:5] <= 3)?
                      3
                    :
                      25
              :
                 (X10[7:4] <= 4)?
                  2
                :
                  1
          :
             (X15[7:6] <= 0)?
               (X6[7:6] <= 3)?
                 (X2[7:6] <= 0)?
                  18
                :
                   (X13[7:6] <= 0)?
                    80
                  :
                     (X2[7:6] <= 1)?
                      3
                    :
                      7
              :
                 (X8[7:5] <= 6)?
                   (X2[7:6] <= 0)?
                    108
                  :
                     (X4[7:6] <= 0)?
                       (X5[7:6] <= 1)?
                        2
                      :
                        16
                    :
                       (X8[7:6] <= 0)?
                         (X0[7:5] <= 0)?
                           (X2[7:5] <= 3)?
                            2
                          :
                            1
                        :
                          46
                      :
                         (X2[7:6] <= 0)?
                          2
                        :
                          3
                :
                   (X2[7:6] <= 0)?
                     (X14[7:6] <= 1)?
                       (X1[7:6] <= 0)?
                        1
                      :
                        8
                    :
                       (X7[7:6] <= 0)?
                        1
                      :
                        4
                  :
                    15
            :
               (X0[7:6] <= 0)?
                27
              :
                1
  :
     (X13[7:5] <= 5)?
       (X0[7:6] <= 0)?
         (X14[7:6] <= 0)?
           (X1[7:4] <= 9)?
             (X8[7:6] <= 2)?
               (X12[7:4] <= 11)?
                34
              :
                 (X5[7:6] <= 2)?
                  1
                :
                  2
            :
              5
          :
             (X3[7:4] <= 13)?
               (X4[7:6] <= 0)?
                2
              :
                8
            :
               (X9[7:6] <= 0)?
                 (X15[7:6] <= 0)?
                  59
                :
                   (X11[7:5] <= 0)?
                    1
                  :
                    1
              :
                2
        :
           (X8[7:5] <= 0)?
             (X0[7:5] <= 0)?
              1
            :
              13
          :
             (X1[7:6] <= 0)?
               (X15[7:6] <= 0)?
                 (X2[7:5] <= 3)?
                  6
                :
                  1
              :
                2
            :
              563
      :
         (X6[7:6] <= 0)?
           (X14[7:6] <= 1)?
             (X9[7:5] <= 1)?
               (X15[7:5] <= 5)?
                324
              :
                1
            :
               (X13[7:5] <= 0)?
                 (X11[7:6] <= 0)?
                  4
                :
                  2
              :
                 (X15[7:6] <= 1)?
                  1
                :
                  12
          :
             (X12[7:5] <= 3)?
              17
            :
              29
        :
           (X15[7:5] <= 1)?
             (X7[7:6] <= 0)?
               (X10[7:6] <= 1)?
                 (X2[7:6] <= 1)?
                  1
                :
                  4
              :
                 (X0[7:6] <= 0)?
                  2
                :
                  3
            :
               (X11[7:6] <= 0)?
                 (X3[7:6] <= 2)?
                   (X4[7:6] <= 0)?
                    1
                  :
                    3
                :
                  4
              :
                6
          :
             (X15[7:6] <= 0)?
               (X7[7:5] <= 0)?
                3
              :
                17
            :
              177
    :
       (X8[7:5] <= 0)?
         (X14[7:6] <= 1)?
           (X12[7:6] <= 0)?
            9
          :
             (X11[7:6] <= 0)?
               (X12[7:5] <= 5)?
                16
              :
                12
            :
               (X1[7:6] <= 0)?
                1
              :
                331
        :
           (X13[7:5] <= 3)?
             (X6[7:5] <= 0)?
              4
            :
               (X11[7:5] <= 1)?
                 (X5[7:6] <= 0)?
                   (X9[7:6] <= 0)?
                    1
                  :
                    1
                :
                  40
              :
                 (X5[7:4] <= 5)?
                  3
                :
                  1
          :
             (X12[7:5] <= 3)?
               (X5[7:5] <= 0)?
                377
              :
                 (X12[7:6] <= 0)?
                  47
                :
                  1
            :
              1
      :
         (X7[7:5] <= 0)?
           (X2[7:6] <= 0)?
             (X6[7:6] <= 4)?
               (X4[7:6] <= 0)?
                716
              :
                 (X3[7:6] <= 1)?
                  1
                :
                  1
            :
               (X15[7:6] <= 3)?
                11
              :
                4
          :
             (X11[7:6] <= 2)?
               (X6[7:6] <= 0)?
                1
              :
                1
            :
              11
        :
           (X9[7:6] <= 0)?
             (X12[7:6] <= 0)?
              1
            :
              31
          :
             (X5[7:5] <= 1)?
               (X6[7:6] <= 0)?
                2
              :
                24
            :
              16
;
endmodule
