module top(X16, out);
input [7:0] X16;
output [3:0] out;
assign out = 
   (X16 <= 14)?
    800
  :
     (X16 <= 43)?
      794
    :
       (X16 <= 71)?
        793
      :
         (X16 <= 185)?
           (X16 <= 128)?
             (X16 <= 100)?
              734
            :
              786
          :
             (X16 <= 156)?
              738
            :
              752
        :
           (X16 <= 213)?
            805
          :
             (X16 <= 242)?
              747
            :
              745
;
endmodule
