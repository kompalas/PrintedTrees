module top(X16, out);
input [7:0] X16;
output [3:0] out;
assign out = 
   (X16[7:5] <= 0)?
    800
  :
     (X16[7:4] <= 0)?
      794
    :
       (X16[7:6] <= 1)?
        793
      :
         (X16[7:4] <= 4)?
           (X16[7:2] <= 48)?
             (X16[7:5] <= 4)?
              734
            :
              786
          :
             (X16[7:6] <= 2)?
              738
            :
              752
        :
           (X16[7:5] <= 6)?
            805
          :
             (X16[7:2] <= 64)?
              747
            :
              745
;
endmodule
