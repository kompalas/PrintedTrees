module top(X0, X1, X2, X3, X4, X5, X6, X7, X8, out);
input [7:0] X0;
input [7:0] X1;
input [7:0] X2;
input [7:0] X3;
input [7:0] X4;
input [7:0] X5;
input [7:0] X6;
input [7:0] X7;
input [7:0] X8;
output [1:0] out;
assign out = 
   (X2[7:6] <= 0)?
     (X6[7:6] <= 1)?
       (X5[7:5] <= 3)?
        291
      :
         (X3[7:6] <= 1)?
          2
        :
          2
    :
       (X7[7:5] <= 1)?
        10
      :
         (X1[7:6] <= 1)?
           (X5[7:6] <= 0)?
             (X3[7:6] <= 1)?
               (X0[7:5] <= 1)?
                5
              :
                 (X6[7:5] <= 3)?
                  3
                :
                   (X4[7:6] <= 3)?
                    3
                  :
                    1
            :
              2
          :
            5
        :
          9
  :
     (X7[7:6] <= 1)?
       (X6[7:6] <= 1)?
         (X1[7:6] <= 3)?
           (X4[7:6] <= 1)?
             (X8[7:6] <= 1)?
               (X3[7:6] <= 1)?
                 (X5[7:5] <= 3)?
                  5
                :
                   (X6[7:4] <= 7)?
                    1
                  :
                    1
              :
                1
            :
              3
          :
            5
        :
          7
      :
        21
    :
      101
;
endmodule
