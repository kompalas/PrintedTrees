module top(X0, X1, X2, X3, X4, X5, out);
input [7:0] X0;
input [7:0] X1;
input [7:0] X2;
input [7:0] X3;
input [7:0] X4;
input [7:0] X5;
output [1:0] out;
assign out = 
   (X5[7:3] <= 2)?
     (X3[7:6] <= 1)?
       (X4[7:3] <= 15)?
        13
      :
         (X1[7:5] <= 3)?
           (X0[7:6] <= 0)?
            1
          :
            11
        :
           (X4[7:5] <= 8)?
             (X1[7:4] <= 8)?
               (X0[7:5] <= 1)?
                 (X5[7:5] <= 0)?
                  8
                :
                   (X4[7:5] <= 3)?
                    1
                  :
                    1
              :
                 (X3[7:4] <= 3)?
                  3
                :
                   (X0[7:5] <= 2)?
                    1
                  :
                    4
            :
              6
          :
             (X5[7:6] <= 1)?
               (X1[7:4] <= 9)?
                7
              :
                1
            :
              2
    :
       (X4[7:5] <= 3)?
         (X3[7:5] <= 3)?
           (X1[7:6] <= 0)?
             (X4[7:6] <= 2)?
              6
            :
               (X5[7:6] <= 1)?
                 (X5[7:4] <= 0)?
                  1
                :
                  3
              :
                3
          :
             (X2[7:5] <= 3)?
              1
            :
              2
        :
           (X0[7:4] <= 9)?
             (X0[7:4] <= 7)?
              2
            :
              2
          :
            5
      :
        29
  :
     (X5[7:4] <= 2)?
       (X5[7:5] <= 2)?
         (X4[7:4] <= 10)?
          24
        :
           (X2[7:5] <= 3)?
            3
          :
            1
      :
        1
    :
      75
;
endmodule
