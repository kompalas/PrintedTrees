module top(X6, X13, X169, X236, X251, X260, X278, out);
input [7:0] X6;
input [7:0] X13;
input [7:0] X169;
input [7:0] X236;
input [7:0] X251;
input [7:0] X260;
input [7:0] X278;
output [4:0] out;
assign out = 
   (X278[7:4] <= -1)?
    165
  :
     (X278[7:5] <= 0)?
      25
    :
       (X278[7:6] <= -1)?
         (X13[7:4] <= -4)?
          19
        :
           (X278[7:5] <= -1)?
            11
          :
             (X169[7:6] <= 0)?
              10
            :
               (X6[7:6] <= -2)?
                10
              :
                 (X236[7:6] <= 0)?
                  4
                :
                   (X251[7:6] <= 0)?
                    2
                  :
                    2
      :
         (X278[7:6] <= -1)?
          31
        :
           (X260[7:5] <= 0)?
            13
          :
            2
;
endmodule
