module top(X6, X13, X169, X236, X251, X260, X278, out);
input [7:0] X6;
input [7:0] X13;
input [7:0] X169;
input [7:0] X236;
input [7:0] X251;
input [7:0] X260;
input [7:0] X278;
output [4:0] out;
assign out = 
   (X278[7:1] <= 2)?
    165
  :
     (X278[7:2] <= 4)?
      25
    :
       (X278[7:2] <= 38)?
         (X13[7:5] <= 3)?
          19
        :
           (X278[7:1] <= 24)?
            11
          :
             (X169[7:4] <= 12)?
              10
            :
               (X6[7:5] <= 2)?
                10
              :
                 (X236[7:4] <= 6)?
                  4
                :
                   (X251 <= 197)?
                    2
                  :
                    2
      :
         (X278[7:6] <= 1)?
          31
        :
           (X260[7:6] <= 6)?
            13
          :
            2
;
endmodule
