module top(X0, X2, X5, X9, X10, X12, X13, X50, X55, X74, X91, X124, X139, X147, X164, X170, X171, X175, X180, X184, X186, X190, X195, X199, X205, X209, X216, X221, X222, X235, X236, X240, X246, X251, X255, X256, X257, X258, X261, X264, X265, X271, X274, X275, X276, out);
input [7:0] X0;
input [7:0] X2;
input [7:0] X5;
input [7:0] X9;
input [7:0] X10;
input [7:0] X12;
input [7:0] X13;
input [7:0] X50;
input [7:0] X55;
input [7:0] X74;
input [7:0] X91;
input [7:0] X124;
input [7:0] X139;
input [7:0] X147;
input [7:0] X164;
input [7:0] X170;
input [7:0] X171;
input [7:0] X175;
input [7:0] X180;
input [7:0] X184;
input [7:0] X186;
input [7:0] X190;
input [7:0] X195;
input [7:0] X199;
input [7:0] X205;
input [7:0] X209;
input [7:0] X216;
input [7:0] X221;
input [7:0] X222;
input [7:0] X235;
input [7:0] X236;
input [7:0] X240;
input [7:0] X246;
input [7:0] X251;
input [7:0] X255;
input [7:0] X256;
input [7:0] X257;
input [7:0] X258;
input [7:0] X261;
input [7:0] X264;
input [7:0] X265;
input [7:0] X271;
input [7:0] X274;
input [7:0] X275;
input [7:0] X276;
output [4:0] out;
assign out = 
   (X195 <= 81)?
     (X13 <= 29)?
       (X264 <= 107)?
         (X240 <= 110)?
          13
        :
          2
      :
        3
    :
       (X222 <= 13)?
         (X246 <= 131)?
           (X0 <= 117)?
             (X2 <= 25)?
               (X124 <= 99)?
                1
              :
                 (X205 <= 75)?
                  1
                :
                  1
            :
              3
          :
             (X164 <= 164)?
               (X170 <= 42)?
                1
              :
                2
            :
               (X199 <= 249)?
                3
              :
                1
        :
           (X13 <= 110)?
             (X235 <= 96)?
               (X221 <= 218)?
                 (X180 <= 54)?
                  1
                :
                  1
              :
                5
            :
               (X74 <= 76)?
                 (X271 <= 242)?
                   (X186 <= 138)?
                     (X221 <= 176)?
                      1
                    :
                      32
                  :
                     (X275 <= 163)?
                       (X175 <= 111)?
                        1
                      :
                        9
                    :
                       (X255 <= 117)?
                        1
                      :
                        4
                :
                   (X5 <= 100)?
                     (X251 <= 247)?
                       (X257 <= 112)?
                        1
                      :
                        88
                    :
                       (X261 <= 253)?
                        2
                      :
                        4
                  :
                     (X274 <= 52)?
                      3
                    :
                       (X139 <= 50)?
                        1
                      :
                        2
              :
                 (X9 <= 111)?
                  3
                :
                   (X170 <= 74)?
                    3
                  :
                    1
          :
             (X184 <= 187)?
              6
            :
               (X171 <= 220)?
                1
              :
                2
      :
         (X12 <= 179)?
           (X2 <= 27)?
            19
          :
            1
        :
           (X271 <= 225)?
            1
          :
             (X91 <= 71)?
              1
            :
              1
  :
     (X236 <= 110)?
       (X50 <= 166)?
         (X147 <= 93)?
          3
        :
          2
      :
        6
    :
       (X209 <= 207)?
         (X255 <= 94)?
          2
        :
           (X216 <= 84)?
            1
          :
            8
      :
         (X190 <= 38)?
           (X0 <= 159)?
             (X10 <= 239)?
              15
            :
              2
          :
             (X265 <= 110)?
               (X216 <= 119)?
                12
              :
                 (X55 <= 6)?
                  4
                :
                  2
            :
              2
        :
           (X258 <= 136)?
             (X5 <= 75)?
              2
            :
              2
          :
             (X276 <= 90)?
              2
            :
               (X256 <= 139)?
                1
              :
                2
;
endmodule
