module top(X0, X2, X5, X9, X10, X12, X13, X50, X55, X74, X91, X124, X139, X147, X164, X170, X171, X175, X180, X184, X186, X190, X195, X199, X205, X209, X216, X221, X222, X235, X236, X240, X246, X251, X255, X256, X257, X258, X261, X264, X265, X271, X274, X275, X276, out);
input [7:0] X0;
input [7:0] X2;
input [7:0] X5;
input [7:0] X9;
input [7:0] X10;
input [7:0] X12;
input [7:0] X13;
input [7:0] X50;
input [7:0] X55;
input [7:0] X74;
input [7:0] X91;
input [7:0] X124;
input [7:0] X139;
input [7:0] X147;
input [7:0] X164;
input [7:0] X170;
input [7:0] X171;
input [7:0] X175;
input [7:0] X180;
input [7:0] X184;
input [7:0] X186;
input [7:0] X190;
input [7:0] X195;
input [7:0] X199;
input [7:0] X205;
input [7:0] X209;
input [7:0] X216;
input [7:0] X221;
input [7:0] X222;
input [7:0] X235;
input [7:0] X236;
input [7:0] X240;
input [7:0] X246;
input [7:0] X251;
input [7:0] X255;
input [7:0] X256;
input [7:0] X257;
input [7:0] X258;
input [7:0] X261;
input [7:0] X264;
input [7:0] X265;
input [7:0] X271;
input [7:0] X274;
input [7:0] X275;
input [7:0] X276;
output [4:0] out;
assign out = 
   (X195[7:6] <= 1)?
     (X13[7:5] <= 0)?
       (X264[7:6] <= 1)?
         (X240[7:5] <= 3)?
          13
        :
          2
      :
        3
    :
       (X222[7:6] <= 0)?
         (X246[7:6] <= 1)?
           (X0[7:5] <= 0)?
             (X2[7:4] <= 0)?
               (X124[7:6] <= 4)?
                1
              :
                 (X205[7:6] <= 0)?
                  1
                :
                  1
            :
              3
          :
             (X164[7:4] <= 7)?
               (X170[7:5] <= 0)?
                1
              :
                2
            :
               (X199[7:6] <= 4)?
                3
              :
                1
        :
           (X13[7:6] <= 0)?
             (X235[7:5] <= 3)?
               (X221[7:5] <= 7)?
                 (X180[7:6] <= 0)?
                  1
                :
                  1
              :
                5
            :
               (X74[7:6] <= 1)?
                 (X271[7:6] <= 1)?
                   (X186[7:6] <= 2)?
                     (X221[7:6] <= 3)?
                      1
                    :
                      32
                  :
                     (X275[7:5] <= 0)?
                       (X175[7:6] <= 1)?
                        1
                      :
                        9
                    :
                       (X255[7:5] <= 2)?
                        1
                      :
                        4
                :
                   (X5[7:6] <= 0)?
                     (X251[7:5] <= 3)?
                       (X257[7:5] <= 3)?
                        1
                      :
                        88
                    :
                       (X261[7:4] <= 16)?
                        2
                      :
                        4
                  :
                     (X274[7:6] <= 0)?
                      3
                    :
                       (X139[7:6] <= 0)?
                        1
                      :
                        2
              :
                 (X9[7:6] <= 0)?
                  3
                :
                   (X170[7:6] <= 0)?
                    3
                  :
                    1
          :
             (X184[7:6] <= 0)?
              6
            :
               (X171[7:5] <= 5)?
                1
              :
                2
      :
         (X12[7:4] <= 11)?
           (X2[7:5] <= 1)?
            19
          :
            1
        :
           (X271[7:6] <= 1)?
            1
          :
             (X91[7:6] <= 1)?
              1
            :
              1
  :
     (X236[7:6] <= 0)?
       (X50[7:6] <= 0)?
         (X147[7:5] <= 3)?
          3
        :
          2
      :
        6
    :
       (X209[7:6] <= 2)?
         (X255[7:6] <= 0)?
          2
        :
           (X216[7:6] <= 1)?
            1
          :
            8
      :
         (X190[7:5] <= 0)?
           (X0[7:6] <= 0)?
             (X10[7:6] <= 3)?
              15
            :
              2
          :
             (X265[7:6] <= 0)?
               (X216[7:6] <= 4)?
                12
              :
                 (X55[7:6] <= 0)?
                  4
                :
                  2
            :
              2
        :
           (X258[7:6] <= 1)?
             (X5[7:4] <= 5)?
              2
            :
              2
          :
             (X276[7:5] <= 0)?
              2
            :
               (X256[7:6] <= 2)?
                1
              :
                2
;
endmodule
