module top(X0, X1, X2, X3, X6, X7, X8, X9, X10, X11, X12, X13, X14, X15, X16, X17, X18, X19, out);
input [7:0] X0;
input [7:0] X1;
input [7:0] X2;
input [7:0] X3;
input [7:0] X6;
input [7:0] X7;
input [7:0] X8;
input [7:0] X9;
input [7:0] X10;
input [7:0] X11;
input [7:0] X12;
input [7:0] X13;
input [7:0] X14;
input [7:0] X15;
input [7:0] X16;
input [7:0] X17;
input [7:0] X18;
input [7:0] X19;
output [1:0] out;
assign out = 
   (X7 <= 163)?
     (X17[7:3] <= 10)?
       (X12[7:2] <= 13)?
         (X8[7:3] <= 31)?
          15
        :
          1
      :
         (X13[7:2] <= 19)?
          1
        :
          3
    :
       (X0[7:4] <= 13)?
         (X6[7:2] <= 6)?
           (X16[7:2] <= 19)?
            1
          :
             (X8[7:3] <= 3)?
               (X16[7:3] <= 22)?
                87
              :
                 (X0[7:2] <= 38)?
                   (X1[7:1] <= 20)?
                     (X17[7:5] <= 6)?
                      1
                    :
                      4
                  :
                    4
                :
                  32
            :
              535
        :
           (X2[7:4] <= 4)?
             (X10[7:3] <= 13)?
              31
            :
               (X14[7:3] <= 4)?
                1
              :
                1
          :
             (X1[7:1] <= 18)?
               (X13[7:4] <= 10)?
                1
              :
                3
            :
               (X19[7:5] <= 2)?
                6
              :
                 (X1[7:4] <= 5)?
                  2
                :
                  1
      :
         (X1[7:3] <= 6)?
           (X18[7:3] <= 23)?
             (X6[7:2] <= 6)?
               (X9[7:1] <= 82)?
                 (X2[7:3] <= 6)?
                  60
                :
                   (X2[7:2] <= 7)?
                    2
                  :
                    1
              :
                2
            :
              4
          :
             (X0[7:3] <= 23)?
               (X3[7:3] <= 17)?
                 (X18[7:2] <= 47)?
                  14
                :
                   (X11[7:2] <= 12)?
                    2
                  :
                    2
              :
                3
            :
               (X9[7:3] <= 23)?
                 (X13 <= 99)?
                   (X3[7:5] <= 1)?
                     (X15[7:3] <= 3)?
                      3
                    :
                       (X16[7:2] <= 54)?
                        1
                      :
                        1
                  :
                    16
                :
                   (X0 <= 231)?
                     (X7[7:3] <= 18)?
                       (X12[7:1] <= 97)?
                        4
                      :
                         (X1[7:3] <= 1)?
                          3
                        :
                          1
                    :
                      6
                  :
                     (X1[7:2] <= 6)?
                      6
                    :
                      1
              :
                4
        :
           (X3[7:3] <= 7)?
             (X9[7:4] <= 1)?
               (X19[7:4] <= 0)?
                2
              :
                33
            :
               (X10[7:4] <= 6)?
                1
              :
                3
          :
             (X15[7:3] <= 2)?
              144
            :
               (X12[7:3] <= 27)?
                5
              :
                1
  :
     (X9[7:2] <= 6)?
       (X17[7:3] <= 10)?
         (X13[7:2] <= 62)?
           (X14[7:4] <= 10)?
            45
          :
             (X6[7:3] <= 7)?
              1
            :
              1
        :
          2
      :
         (X7[7:2] <= 56)?
           (X19[7:2] <= 1)?
             (X12[7:4] <= 5)?
              5
            :
               (X3[7:3] <= 7)?
                 (X7 <= 185)?
                  2
                :
                  4
              :
                22
          :
             (X6[7:1] <= 39)?
              112
            :
               (X2[7:3] <= 4)?
                3
              :
                2
        :
           (X18[7:5] <= 8)?
            5
          :
            3
    :
       (X9[7:2] <= 48)?
         (X7[7:2] <= 58)?
           (X0[7:4] <= 11)?
             (X8[7:1] <= 7)?
               (X3[7:2] <= 23)?
                 (X1[7:1] <= 19)?
                   (X7[7:4] <= 16)?
                    26
                  :
                     (X9[7:3] <= 15)?
                      1
                    :
                      1
                :
                  2
              :
                 (X14 <= 114)?
                  4
                :
                  1
            :
               (X14[7:5] <= 5)?
                16
              :
                2
          :
             (X9[7:4] <= 2)?
               (X7 <= 192)?
                 (X9[7:3] <= 10)?
                   (X16[7:5] <= 8)?
                    37
                  :
                     (X1[7:2] <= 2)?
                      2
                    :
                      1
                :
                  1
              :
                 (X13[7:2] <= 24)?
                   (X2[7:3] <= 2)?
                    4
                  :
                    3
                :
                  4
            :
              82
        :
           (X3[7:1] <= 26)?
            8
          :
            2
      :
         (X3[7:3] <= 14)?
          24
        :
           (X8[7:4] <= 3)?
            1
          :
            2
;
endmodule
