module top(X0, X1, X4, X9, X12, X28, X30, X32, X37, X38, X41, X42, X44, X49, X51, X52, X54, X55, X56, X57, X58, X62, X63, X65, X69, X73, X90, X93, X101, X102, X106, X113, X114, X115, X118, X125, X128, X133, X136, X137, X139, X141, X142, X147, X148, X155, X159, X161, X162, X165, X169, X170, X172, X180, X181, X185, X190, X192, X198, X199, X209, X210, X227, X238, X240, X244, X245, X248, X258, X259, X263, X265, X268, X270, X273, X274, X275, X276, X283, X286, X287, X290, X296, X300, X301, X302, X310, X312, X313, X319, X320, X323, X324, X326, X327, X330, X331, X335, X336, X340, X342, X358, X361, X362, X370, X371, X376, X380, X387, X388, X394, X395, X403, X405, X409, X410, X414, X428, X432, X434, X435, X445, X449, X452, X455, X457, X458, X460, X462, X477, X481, X483, X488, X489, X498, X504, X509, X514, X524, X527, X535, X537, X539, X542, X550, X554, X558, X560, out);
input [7:0] X0;
input [7:0] X1;
input [7:0] X4;
input [7:0] X9;
input [7:0] X12;
input [7:0] X28;
input [7:0] X30;
input [7:0] X32;
input [7:0] X37;
input [7:0] X38;
input [7:0] X41;
input [7:0] X42;
input [7:0] X44;
input [7:0] X49;
input [7:0] X51;
input [7:0] X52;
input [7:0] X54;
input [7:0] X55;
input [7:0] X56;
input [7:0] X57;
input [7:0] X58;
input [7:0] X62;
input [7:0] X63;
input [7:0] X65;
input [7:0] X69;
input [7:0] X73;
input [7:0] X90;
input [7:0] X93;
input [7:0] X101;
input [7:0] X102;
input [7:0] X106;
input [7:0] X113;
input [7:0] X114;
input [7:0] X115;
input [7:0] X118;
input [7:0] X125;
input [7:0] X128;
input [7:0] X133;
input [7:0] X136;
input [7:0] X137;
input [7:0] X139;
input [7:0] X141;
input [7:0] X142;
input [7:0] X147;
input [7:0] X148;
input [7:0] X155;
input [7:0] X159;
input [7:0] X161;
input [7:0] X162;
input [7:0] X165;
input [7:0] X169;
input [7:0] X170;
input [7:0] X172;
input [7:0] X180;
input [7:0] X181;
input [7:0] X185;
input [7:0] X190;
input [7:0] X192;
input [7:0] X198;
input [7:0] X199;
input [7:0] X209;
input [7:0] X210;
input [7:0] X227;
input [7:0] X238;
input [7:0] X240;
input [7:0] X244;
input [7:0] X245;
input [7:0] X248;
input [7:0] X258;
input [7:0] X259;
input [7:0] X263;
input [7:0] X265;
input [7:0] X268;
input [7:0] X270;
input [7:0] X273;
input [7:0] X274;
input [7:0] X275;
input [7:0] X276;
input [7:0] X283;
input [7:0] X286;
input [7:0] X287;
input [7:0] X290;
input [7:0] X296;
input [7:0] X300;
input [7:0] X301;
input [7:0] X302;
input [7:0] X310;
input [7:0] X312;
input [7:0] X313;
input [7:0] X319;
input [7:0] X320;
input [7:0] X323;
input [7:0] X324;
input [7:0] X326;
input [7:0] X327;
input [7:0] X330;
input [7:0] X331;
input [7:0] X335;
input [7:0] X336;
input [7:0] X340;
input [7:0] X342;
input [7:0] X358;
input [7:0] X361;
input [7:0] X362;
input [7:0] X370;
input [7:0] X371;
input [7:0] X376;
input [7:0] X380;
input [7:0] X387;
input [7:0] X388;
input [7:0] X394;
input [7:0] X395;
input [7:0] X403;
input [7:0] X405;
input [7:0] X409;
input [7:0] X410;
input [7:0] X414;
input [7:0] X428;
input [7:0] X432;
input [7:0] X434;
input [7:0] X435;
input [7:0] X445;
input [7:0] X449;
input [7:0] X452;
input [7:0] X455;
input [7:0] X457;
input [7:0] X458;
input [7:0] X460;
input [7:0] X462;
input [7:0] X477;
input [7:0] X481;
input [7:0] X483;
input [7:0] X488;
input [7:0] X489;
input [7:0] X498;
input [7:0] X504;
input [7:0] X509;
input [7:0] X514;
input [7:0] X524;
input [7:0] X527;
input [7:0] X535;
input [7:0] X537;
input [7:0] X539;
input [7:0] X542;
input [7:0] X550;
input [7:0] X554;
input [7:0] X558;
input [7:0] X560;
output [2:0] out;
assign out = 
   (X102 <= 157)?
     (X56 <= 89)?
       (X63 <= 62)?
         (X118 <= 203)?
           (X137 <= 7)?
             (X301 <= 3)?
               (X310 <= 0)?
                8
              :
                1
            :
              335
          :
            1
        :
           (X327 <= 2)?
             (X210 <= 133)?
              3
            :
              1
          :
            5
      :
         (X58 <= 138)?
           (X51 <= 198)?
             (X113 <= 145)?
              17
            :
              1
          :
             (X198 <= 100)?
              3
            :
              19
        :
           (X560 <= 21)?
            6
          :
             (X106 <= 92)?
              1
            :
              22
    :
       (X560 <= 147)?
         (X49 <= 219)?
          184
        :
           (X340 <= 0)?
             (X445 <= 28)?
              6
            :
               (X199 <= 194)?
                24
              :
                3
          :
             (X481 <= 1)?
               (X63 <= 68)?
                92
              :
                 (X312 <= 0)?
                  4
                :
                  9
            :
               (X32 <= 147)?
                 (X326 <= 16)?
                  2
                :
                  2
              :
                2
      :
         (X139 <= 1)?
           (X58 <= 6)?
             (X403 <= 0)?
               (X57 <= 3)?
                 (X361 <= 0)?
                  11
                :
                  1
              :
                 (X259 <= 2)?
                  10
                :
                  1
            :
               (X320 <= 0)?
                80
              :
                 (X286 <= 2)?
                  6
                :
                   (X118 <= 108)?
                     (X300 <= 141)?
                      3
                    :
                      3
                  :
                    29
          :
             (X41 <= 114)?
              6
            :
               (X142 <= 27)?
                2
              :
                30
        :
           (X51 <= 105)?
             (X245 <= 9)?
               (X42 <= 32)?
                9
              :
                 (X41 <= 138)?
                   (X460 <= 0)?
                     (X125 <= 1)?
                      12
                    :
                       (X394 <= 0)?
                        10
                      :
                        2
                  :
                     (X65 <= 48)?
                       (X558 <= 16)?
                        6
                      :
                         (X263 <= 152)?
                          36
                        :
                           (X380 <= 25)?
                            3
                          :
                            1
                    :
                       (X527 <= 72)?
                        232
                      :
                         (X388 <= 0)?
                           (X319 <= 0)?
                            1
                          :
                            33
                        :
                          2
                :
                   (X57 <= 13)?
                     (X192 <= 159)?
                      23
                    :
                      4
                  :
                     (X539 <= 154)?
                      44
                    :
                      3
            :
               (X488 <= 2)?
                2
              :
                 (X93 <= 212)?
                  1
                :
                  1
          :
             (X248 <= 90)?
               (X498 <= 0)?
                 (X414 <= 0)?
                  37
                :
                  1
              :
                 (X275 <= 31)?
                  7
                :
                  4
            :
               (X101 <= 25)?
                 (X54 <= 121)?
                   (X290 <= 35)?
                     (X161 <= 87)?
                      5
                    :
                       (X190 <= 157)?
                        14
                      :
                        2
                  :
                    13
                :
                   (X335 <= 0)?
                    46
                  :
                     (X169 <= 3)?
                      5
                    :
                      7
              :
                 (X376 <= 6)?
                  2
                :
                  2
  :
     (X69 <= 66)?
       (X302 <= 5)?
         (X38 <= 125)?
           (X395 <= 14)?
             (X268 <= 32)?
              5
            :
              10
          :
             (X30 <= 143)?
               (X537 <= 6)?
                2
              :
                1
            :
              7
        :
           (X455 <= 190)?
            37
          :
            1
      :
         (X52 <= 172)?
           (X159 <= 95)?
             (X371 <= 91)?
              5
            :
               (X358 <= 57)?
                10
              :
                3
          :
             (X457 <= 19)?
               (X41 <= 135)?
                2
              :
                5
            :
               (X136 <= 29)?
                 (X240 <= 25)?
                   (X273 <= 144)?
                    1
                  :
                    1
                :
                  16
              :
                 (X313 <= 3)?
                  1
                :
                  3
        :
           (X434 <= 29)?
             (X73 <= 61)?
               (X449 <= 28)?
                 (X287 <= 207)?
                   (X524 <= 4)?
                    1
                  :
                    23
                :
                  3
              :
                 (X0 <= 153)?
                  10
                :
                  2
            :
              30
          :
             (X37 <= 199)?
               (X457 <= 35)?
                 (X128 <= 49)?
                   (X462 <= 13)?
                    7
                  :
                    3
                :
                   (X192 <= 103)?
                     (X244 <= 88)?
                      6
                    :
                      3
                  :
                    59
              :
                113
            :
               (X403 <= 11)?
                1
              :
                9
    :
       (X509 <= 76)?
         (X37 <= 163)?
           (X69 <= 98)?
             (X394 <= 9)?
               (X265 <= 70)?
                 (X90 <= 43)?
                   (X336 <= 6)?
                    2
                  :
                     (X4 <= 53)?
                      1
                    :
                      2
                :
                  50
              :
                 (X54 <= 92)?
                  12
                :
                   (X49 <= 235)?
                    8
                  :
                    2
            :
               (X57 <= 3)?
                 (X209 <= 174)?
                   (X12 <= 143)?
                    9
                  :
                     (X312 <= 12)?
                      4
                    :
                       (X62 <= 119)?
                        16
                      :
                        2
                :
                   (X428 <= 21)?
                    1
                  :
                    34
              :
                 (X283 <= 14)?
                   (X483 <= 7)?
                     (X1 <= 123)?
                      4
                    :
                       (X324 <= 40)?
                        31
                      :
                        1
                  :
                     (X504 <= 72)?
                      12
                    :
                       (X550 <= 14)?
                        3
                      :
                        1
                :
                   (X342 <= 22)?
                     (X181 <= 90)?
                       (X55 <= 173)?
                         (X435 <= 24)?
                           (X535 <= 76)?
                            8
                          :
                            1
                        :
                           (X258 <= 31)?
                            5
                          :
                            3
                      :
                        19
                    :
                       (X1 <= 123)?
                        2
                      :
                        12
                  :
                    31
          :
             (X44 <= 8)?
               (X488 <= 2)?
                 (X331 <= 29)?
                  4
                :
                   (X133 <= 221)?
                    2
                  :
                     (X57 <= 21)?
                      1
                    :
                      1
              :
                 (X274 <= 90)?
                   (X162 <= 188)?
                    189
                  :
                     (X147 <= 159)?
                       (X185 <= 186)?
                        22
                      :
                        1
                    :
                      2
                :
                  2
            :
               (X181 <= 103)?
                 (X452 <= 117)?
                   (X276 <= 39)?
                     (X90 <= 73)?
                      5
                    :
                       (X165 <= 45)?
                         (X477 <= 16)?
                          3
                        :
                          1
                      :
                        10
                  :
                     (X405 <= 15)?
                       (X409 <= 61)?
                        8
                      :
                        2
                    :
                      9
                :
                   (X28 <= 185)?
                     (X141 <= 29)?
                      1
                    :
                      23
                  :
                    2
              :
                 (X180 <= 139)?
                  44
                :
                  2
        :
           (X409 <= 27)?
             (X296 <= 41)?
               (X452 <= 157)?
                1
              :
                1
            :
              57
          :
             (X159 <= 161)?
               (X199 <= 144)?
                 (X238 <= 168)?
                  21
                :
                   (X410 <= 28)?
                     (X115 <= 130)?
                      3
                    :
                      2
                  :
                     (X458 <= 77)?
                      1
                    :
                      7
              :
                 (X550 <= 4)?
                  1
                :
                  13
            :
               (X170 <= 16)?
                 (X387 <= 5)?
                  2
                :
                  1
              :
                 (X102 <= 231)?
                  24
                :
                  1
      :
         (X57 <= 10)?
           (X514 <= 76)?
             (X9 <= 91)?
               (X172 <= 213)?
                 (X227 <= 140)?
                  16
                :
                  3
              :
                 (X155 <= 79)?
                  1
                :
                  6
            :
               (X115 <= 145)?
                 (X114 <= 50)?
                  1
                :
                  136
              :
                 (X542 <= 63)?
                  3
                :
                  2
          :
             (X432 <= 56)?
               (X170 <= 41)?
                3
              :
                1
            :
               (X458 <= 78)?
                1
              :
                20
        :
           (X330 <= 8)?
             (X489 <= 23)?
              48
            :
              1
          :
             (X38 <= 75)?
               (X238 <= 156)?
                 (X199 <= 129)?
                  32
                :
                  3
              :
                 (X554 <= 157)?
                  9
                :
                  2
            :
               (X270 <= 68)?
                 (X434 <= 37)?
                   (X185 <= 144)?
                     (X323 <= 1)?
                      2
                    :
                      8
                  :
                     (X148 <= 69)?
                      1
                    :
                      6
                :
                   (X370 <= 95)?
                    12
                  :
                    3
              :
                 (X362 <= 215)?
                  27
                :
                  1
;
endmodule
