module top(X6, X13, X169, X236, X251, X260, X278, out);
input [7:0] X6;
input [7:0] X13;
input [7:0] X169;
input [7:0] X236;
input [7:0] X251;
input [7:0] X260;
input [7:0] X278;
output [4:0] out;
assign out = 
   (X278 <= 9)?
    165
  :
     (X278 <= 26)?
      25
    :
       (X278 <= 145)?
         (X13 <= 33)?
          19
        :
           (X278 <= 43)?
            11
          :
             (X169 <= 184)?
              10
            :
               (X6 <= 113)?
                10
              :
                 (X236 <= 115)?
                  4
                :
                   (X251 <= 199)?
                    2
                  :
                    2
      :
         (X278 <= 188)?
          31
        :
           (X260 <= 179)?
            13
          :
            2
;
endmodule
