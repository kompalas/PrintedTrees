module top(X2, X6, X9, X10, X12, X14, X23, X28, X32, X36, X37, X40, X41, X42, X43, X50, X51, X54, X55, X56, X57, X58, X63, X65, X68, X69, X74, X76, X77, X86, X88, X89, X100, X102, X111, X115, X117, X118, X128, X131, X133, X139, X140, X141, X144, X145, X147, X150, X152, X158, X175, X178, X179, X181, X185, X187, X189, X196, X197, X198, X203, X204, X214, X221, X224, X230, X238, X243, X246, X252, X257, X264, X266, X270, X276, X280, X288, X293, X295, X300, X301, X302, X305, X306, X317, X321, X330, X331, X335, X339, X343, X357, X358, X365, X369, X371, X374, X387, X390, X394, X396, X407, X410, X415, X417, X418, X427, X434, X435, X440, X448, X449, X453, X454, X464, X467, X476, X485, X486, X490, X491, X492, X494, X498, X504, X507, X509, X510, X515, X536, X546, X552, X554, X555, X557, X558, X559, X560, out);
input [7:0] X2;
input [7:0] X6;
input [7:0] X9;
input [7:0] X10;
input [7:0] X12;
input [7:0] X14;
input [7:0] X23;
input [7:0] X28;
input [7:0] X32;
input [7:0] X36;
input [7:0] X37;
input [7:0] X40;
input [7:0] X41;
input [7:0] X42;
input [7:0] X43;
input [7:0] X50;
input [7:0] X51;
input [7:0] X54;
input [7:0] X55;
input [7:0] X56;
input [7:0] X57;
input [7:0] X58;
input [7:0] X63;
input [7:0] X65;
input [7:0] X68;
input [7:0] X69;
input [7:0] X74;
input [7:0] X76;
input [7:0] X77;
input [7:0] X86;
input [7:0] X88;
input [7:0] X89;
input [7:0] X100;
input [7:0] X102;
input [7:0] X111;
input [7:0] X115;
input [7:0] X117;
input [7:0] X118;
input [7:0] X128;
input [7:0] X131;
input [7:0] X133;
input [7:0] X139;
input [7:0] X140;
input [7:0] X141;
input [7:0] X144;
input [7:0] X145;
input [7:0] X147;
input [7:0] X150;
input [7:0] X152;
input [7:0] X158;
input [7:0] X175;
input [7:0] X178;
input [7:0] X179;
input [7:0] X181;
input [7:0] X185;
input [7:0] X187;
input [7:0] X189;
input [7:0] X196;
input [7:0] X197;
input [7:0] X198;
input [7:0] X203;
input [7:0] X204;
input [7:0] X214;
input [7:0] X221;
input [7:0] X224;
input [7:0] X230;
input [7:0] X238;
input [7:0] X243;
input [7:0] X246;
input [7:0] X252;
input [7:0] X257;
input [7:0] X264;
input [7:0] X266;
input [7:0] X270;
input [7:0] X276;
input [7:0] X280;
input [7:0] X288;
input [7:0] X293;
input [7:0] X295;
input [7:0] X300;
input [7:0] X301;
input [7:0] X302;
input [7:0] X305;
input [7:0] X306;
input [7:0] X317;
input [7:0] X321;
input [7:0] X330;
input [7:0] X331;
input [7:0] X335;
input [7:0] X339;
input [7:0] X343;
input [7:0] X357;
input [7:0] X358;
input [7:0] X365;
input [7:0] X369;
input [7:0] X371;
input [7:0] X374;
input [7:0] X387;
input [7:0] X390;
input [7:0] X394;
input [7:0] X396;
input [7:0] X407;
input [7:0] X410;
input [7:0] X415;
input [7:0] X417;
input [7:0] X418;
input [7:0] X427;
input [7:0] X434;
input [7:0] X435;
input [7:0] X440;
input [7:0] X448;
input [7:0] X449;
input [7:0] X453;
input [7:0] X454;
input [7:0] X464;
input [7:0] X467;
input [7:0] X476;
input [7:0] X485;
input [7:0] X486;
input [7:0] X490;
input [7:0] X491;
input [7:0] X492;
input [7:0] X494;
input [7:0] X498;
input [7:0] X504;
input [7:0] X507;
input [7:0] X509;
input [7:0] X510;
input [7:0] X515;
input [7:0] X536;
input [7:0] X546;
input [7:0] X552;
input [7:0] X554;
input [7:0] X555;
input [7:0] X557;
input [7:0] X558;
input [7:0] X559;
input [7:0] X560;
output [2:0] out;
assign out = 
   (X102 <= 158)?
     (X56 <= 70)?
       (X63 <= 61)?
         (X118 <= 203)?
           (X88 <= 86)?
            336
          :
            1
        :
           (X293 <= 118)?
            3
          :
            3
      :
         (X54 <= 227)?
           (X51 <= 196)?
            16
          :
             (X198 <= 100)?
              4
            :
              24
        :
           (X55 <= 147)?
            7
          :
            25
    :
       (X51 <= 130)?
         (X139 <= 1)?
           (X58 <= 6)?
             (X139 <= 0)?
              53
            :
               (X417 <= 0)?
                 (X57 <= 4)?
                   (X453 <= 138)?
                    28
                  :
                     (X252 <= 1)?
                      8
                    :
                      3
                :
                   (X306 <= 0)?
                    15
                  :
                    2
              :
                 (X14 <= 237)?
                   (X305 <= 0)?
                    3
                  :
                    2
                :
                  54
          :
             (X41 <= 114)?
              14
            :
              29
        :
           (X181 <= 20)?
             (X51 <= 106)?
               (X54 <= 32)?
                11
              :
                 (X50 <= 138)?
                   (X448 <= 52)?
                     (X435 <= 0)?
                       (X147 <= 136)?
                         (X536 <= 152)?
                          32
                        :
                          1
                      :
                         (X554 <= 132)?
                          6
                        :
                          3
                    :
                       (X115 <= 85)?
                         (X144 <= 90)?
                           (X357 <= 2)?
                            3
                          :
                            4
                        :
                          26
                      :
                        256
                  :
                     (X115 <= 115)?
                       (X485 <= 0)?
                        8
                      :
                        2
                    :
                      8
                :
                   (X559 <= 116)?
                     (X187 <= 45)?
                      1
                    :
                      37
                  :
                     (X54 <= 78)?
                       (X23 <= 45)?
                        2
                      :
                        8
                    :
                       (X434 <= 15)?
                        24
                      :
                        1
            :
               (X560 <= 161)?
                 (X40 <= 249)?
                   (X32 <= 150)?
                    45
                  :
                     (X14 <= 240)?
                       (X557 <= 33)?
                        1
                      :
                        4
                    :
                      8
                :
                  10
              :
                 (X189 <= 94)?
                   (X492 <= 0)?
                    1
                  :
                    35
                :
                   (X224 <= 106)?
                    6
                  :
                     (X300 <= 80)?
                       (X554 <= 196)?
                        3
                      :
                        1
                    :
                      13
          :
             (X150 <= 161)?
               (X498 <= 3)?
                3
              :
                4
            :
               (X196 <= 113)?
                 (X214 <= 110)?
                  3
                :
                  1
              :
                6
      :
         (X57 <= 5)?
           (X41 <= 100)?
            18
          :
             (X145 <= 148)?
               (X41 <= 123)?
                7
              :
                8
            :
              54
        :
           (X179 <= 22)?
             (X36 <= 51)?
               (X214 <= 7)?
                3
              :
                2
            :
              232
          :
             (X427 <= 45)?
              2
            :
              3
  :
     (X65 <= 75)?
       (X69 <= 62)?
         (X560 <= 132)?
           (X371 <= 91)?
             (X264 <= 105)?
              2
            :
              5
          :
             (X494 <= 5)?
              10
            :
               (X65 <= 28)?
                2
              :
                2
        :
           (X330 <= 6)?
             (X490 <= 7)?
              18
            :
               (X507 <= 52)?
                1
              :
                3
          :
             (X158 <= 155)?
               (X246 <= 85)?
                 (X515 <= 143)?
                  109
                :
                  1
              :
                 (X203 <= 73)?
                  2
                :
                   (X407 <= 31)?
                    1
                  :
                    1
            :
               (X486 <= 11)?
                 (X12 <= 189)?
                   (X89 <= 61)?
                     (X491 <= 24)?
                      12
                    :
                      1
                  :
                     (X302 <= 86)?
                      10
                    :
                      1
                :
                   (X331 <= 18)?
                    1
                  :
                    4
              :
                25
      :
         (X330 <= 10)?
           (X434 <= 43)?
             (X28 <= 123)?
               (X343 <= 12)?
                2
              :
                 (X270 <= 46)?
                  2
                :
                  2
            :
               (X77 <= 255)?
                103
              :
                1
          :
             (X276 <= 28)?
              7
            :
               (X185 <= 175)?
                10
              :
                1
        :
           (X57 <= 4)?
             (X257 <= 168)?
               (X464 <= 10)?
                 (X175 <= 79)?
                   (X74 <= 200)?
                    4
                  :
                    2
                :
                   (X288 <= 219)?
                    8
                  :
                    1
              :
                 (X390 <= 14)?
                  1
                :
                  31
            :
               (X335 <= 20)?
                2
              :
                21
          :
             (X14 <= 115)?
               (X374 <= 64)?
                5
              :
                34
            :
               (X40 <= 207)?
                 (X76 <= 182)?
                  3
                :
                   (X140 <= 76)?
                    14
                  :
                    2
              :
                 (X203 <= 61)?
                   (X41 <= 148)?
                    3
                  :
                    10
                :
                   (X552 <= 147)?
                     (X238 <= 135)?
                       (X295 <= 87)?
                         (X141 <= 40)?
                          1
                        :
                          20
                      :
                         (X230 <= 64)?
                           (X117 <= 80)?
                            1
                          :
                            8
                        :
                          6
                    :
                       (X56 <= 237)?
                        72
                      :
                        1
                  :
                     (X243 <= 71)?
                      1
                    :
                      4
    :
       (X509 <= 81)?
         (X37 <= 163)?
           (X476 <= 5)?
             (X394 <= 10)?
               (X102 <= 216)?
                 (X560 <= 153)?
                  3
                :
                   (X221 <= 203)?
                     (X339 <= 14)?
                      4
                    :
                      4
                  :
                    57
              :
                3
            :
               (X317 <= 22)?
                 (X449 <= 20)?
                   (X387 <= 3)?
                    2
                  :
                    39
                :
                   (X102 <= 209)?
                    8
                  :
                     (X396 <= 8)?
                      1
                    :
                      2
              :
                 (X427 <= 40)?
                   (X100 <= 87)?
                    24
                  :
                     (X369 <= 74)?
                       (X152 <= 137)?
                        2
                      :
                        7
                    :
                      13
                :
                   (X178 <= 7)?
                     (X358 <= 3)?
                      1
                    :
                      8
                  :
                     (X204 <= 22)?
                       (X266 <= 110)?
                        3
                      :
                        1
                    :
                       (X128 <= 44)?
                         (X546 <= 39)?
                          1
                        :
                          2
                      :
                        17
          :
             (X41 <= 78)?
              13
            :
               (X42 <= 133)?
                 (X559 <= 121)?
                   (X43 <= 5)?
                     (X440 <= 32)?
                       (X10 <= 65)?
                         (X510 <= 175)?
                          4
                        :
                          3
                      :
                        69
                    :
                      3
                  :
                     (X28 <= 157)?
                       (X68 <= 204)?
                         (X418 <= 56)?
                          11
                        :
                          2
                      :
                        4
                    :
                       (X280 <= 101)?
                        3
                      :
                        7
                :
                   (X434 <= 26)?
                     (X6 <= 77)?
                       (X133 <= 207)?
                         (X558 <= 41)?
                          3
                        :
                          1
                      :
                        46
                    :
                      7
                  :
                     (X467 <= 0)?
                       (X68 <= 198)?
                        4
                      :
                        2
                    :
                       (X555 <= 28)?
                         (X2 <= 79)?
                          2
                        :
                          9
                      :
                        192
              :
                 (X111 <= 152)?
                  5
                :
                  5
        :
           (X55 <= 175)?
             (X197 <= 113)?
               (X41 <= 105)?
                 (X415 <= 11)?
                  1
                :
                  1
              :
                23
            :
               (X2 <= 82)?
                4
              :
                 (X50 <= 166)?
                  20
                :
                   (X86 <= 88)?
                    1
                  :
                    1
          :
             (X41 <= 170)?
               (X158 <= 195)?
                27
              :
                 (X454 <= 108)?
                  1
                :
                  1
            :
              17
      :
         (X9 <= 124)?
           (X50 <= 84)?
            9
          :
             (X276 <= 59)?
               (X321 <= 34)?
                 (X560 <= 207)?
                  32
                :
                  2
              :
                 (X504 <= 95)?
                   (X410 <= 65)?
                     (X365 <= 95)?
                      3
                    :
                      13
                  :
                     (X301 <= 8)?
                      1
                    :
                      5
                :
                  13
            :
               (X131 <= 26)?
                1
              :
                7
        :
          66
;
endmodule
