module top(X0, X1, X2, X3, X4, out);
input [7:0] X0;
input [7:0] X1;
input [7:0] X2;
input [7:0] X3;
input [7:0] X4;
output [0:0] out;
assign out = 
   (X0 <= 21)?
     (X2 <= 128)?
       (X1 <= 153)?
         (X3 <= 160)?
           (X4 <= 43)?
            1
          :
             (X1 <= 54)?
              42
            :
               (X1 <= 133)?
                 (X4 <= 128)?
                  17
                :
                   (X1 <= 130)?
                     (X1 <= 84)?
                       (X1 <= 74)?
                         (X1 <= 57)?
                           (X2 <= 43)?
                            3
                          :
                            2
                        :
                          17
                      :
                         (X0 <= 16)?
                          3
                        :
                           (X3 <= 32)?
                             (X1 <= 77)?
                               (X2 <= 43)?
                                3
                              :
                                4
                            :
                               (X2 <= 43)?
                                 (X1 <= 80)?
                                  2
                                :
                                  3
                              :
                                2
                          :
                            2
                    :
                       (X1 <= 113)?
                        40
                      :
                         (X1 <= 120)?
                           (X2 <= 43)?
                             (X1 <= 117)?
                              1
                            :
                              6
                          :
                            4
                        :
                          12
                  :
                     (X2 <= 43)?
                      2
                    :
                      1
              :
                22
        :
           (X1 <= 121)?
            5
          :
             (X3 <= 224)?
               (X2 <= 43)?
                1
              :
                 (X1 <= 131)?
                   (X1 <= 126)?
                    1
                  :
                    2
                :
                   (X1 <= 148)?
                     (X1 <= 139)?
                      1
                    :
                      1
                  :
                    2
            :
              1
      :
         (X1 <= 176)?
           (X1 <= 172)?
             (X2 <= 43)?
               (X4 <= 85)?
                1
              :
                 (X3 <= 128)?
                   (X3 <= 32)?
                     (X1 <= 166)?
                       (X1 <= 156)?
                        1
                      :
                         (X0 <= 16)?
                          1
                        :
                           (X1 <= 161)?
                            1
                          :
                            2
                    :
                      1
                  :
                    1
                :
                  1
            :
               (X3 <= 160)?
                5
              :
                1
          :
            2
        :
           (X4 <= 43)?
             (X1 <= 190)?
              1
            :
              1
          :
            9
    :
       (X1 <= 159)?
         (X1 <= 123)?
           (X1 <= 113)?
             (X1 <= 31)?
              2
            :
               (X1 <= 39)?
                1
              :
                 (X1 <= 110)?
                   (X1 <= 100)?
                     (X1 <= 74)?
                       (X3 <= 224)?
                        6
                      :
                        1
                    :
                       (X0 <= 12)?
                        1
                      :
                         (X3 <= 224)?
                           (X1 <= 97)?
                             (X3 <= 160)?
                               (X3 <= 64)?
                                 (X1 <= 85)?
                                  2
                                :
                                  2
                              :
                                 (X1 <= 87)?
                                  2
                                :
                                  1
                            :
                               (X1 <= 84)?
                                 (X4 <= 128)?
                                  1
                                :
                                  1
                              :
                                3
                          :
                            2
                        :
                          1
                  :
                     (X3 <= 224)?
                      6
                    :
                      1
                :
                   (X2 <= 213)?
                    1
                  :
                    2
          :
            6
        :
           (X1 <= 156)?
             (X1 <= 130)?
               (X4 <= 213)?
                 (X1 <= 126)?
                  1
                :
                   (X2 <= 213)?
                    1
                  :
                     (X3 <= 160)?
                      1
                    :
                      1
              :
                1
            :
               (X1 <= 139)?
                 (X3 <= 160)?
                  3
                :
                   (X1 <= 133)?
                    1
                  :
                     (X3 <= 224)?
                       (X2 <= 213)?
                        1
                      :
                        1
                    :
                      2
              :
                 (X3 <= 64)?
                  1
                :
                   (X4 <= 128)?
                    1
                  :
                     (X0 <= 16)?
                      1
                    :
                       (X3 <= 224)?
                         (X1 <= 149)?
                           (X3 <= 160)?
                            2
                          :
                             (X1 <= 146)?
                               (X2 <= 213)?
                                1
                              :
                                1
                            :
                              2
                        :
                           (X2 <= 213)?
                            2
                          :
                             (X1 <= 153)?
                               (X3 <= 160)?
                                1
                              :
                                1
                            :
                              1
                      :
                         (X1 <= 148)?
                          1
                        :
                          2
          :
            3
      :
         (X1 <= 192)?
           (X0 <= 9)?
            3
          :
             (X1 <= 179)?
               (X1 <= 169)?
                 (X1 <= 166)?
                   (X3 <= 96)?
                    1
                  :
                     (X1 <= 162)?
                       (X3 <= 224)?
                        2
                      :
                        1
                    :
                       (X3 <= 224)?
                        2
                      :
                        1
                :
                  1
              :
                6
            :
               (X4 <= 128)?
                1
              :
                 (X3 <= 32)?
                  1
                :
                   (X3 <= 96)?
                    1
                  :
                     (X2 <= 213)?
                      1
                    :
                       (X3 <= 160)?
                         (X1 <= 185)?
                          1
                        :
                          1
                      :
                        1
        :
          4
  :
     (X4 <= 213)?
       (X3 <= 32)?
         (X0 <= 26)?
           (X2 <= 128)?
            5
          :
             (X4 <= 85)?
              1
            :
              1
        :
          2
      :
         (X1 <= 56)?
           (X2 <= 171)?
            1
          :
            1
        :
           (X4 <= 128)?
             (X2 <= 128)?
              1
            :
               (X1 <= 139)?
                 (X1 <= 130)?
                  3
                :
                  1
              :
                4
          :
             (X1 <= 215)?
               (X1 <= 179)?
                 (X1 <= 113)?
                   (X1 <= 80)?
                     (X1 <= 75)?
                      5
                    :
                       (X3 <= 224)?
                        1
                      :
                        1
                  :
                    27
                :
                   (X1 <= 120)?
                     (X2 <= 213)?
                      1
                    :
                       (X1 <= 117)?
                         (X3 <= 192)?
                          1
                        :
                          1
                      :
                         (X3 <= 160)?
                          1
                        :
                          3
                  :
                     (X1 <= 123)?
                      10
                    :
                       (X1 <= 126)?
                         (X2 <= 171)?
                          1
                        :
                          1
                      :
                         (X3 <= 96)?
                           (X1 <= 148)?
                            1
                          :
                            3
                        :
                           (X1 <= 143)?
                            19
                          :
                             (X3 <= 160)?
                              15
                            :
                               (X1 <= 176)?
                                 (X1 <= 159)?
                                   (X1 <= 146)?
                                     (X3 <= 224)?
                                      1
                                    :
                                      2
                                  :
                                     (X1 <= 153)?
                                      6
                                    :
                                       (X3 <= 224)?
                                         (X1 <= 156)?
                                          2
                                        :
                                          6
                                      :
                                         (X1 <= 156)?
                                          3
                                        :
                                          1
                                :
                                   (X1 <= 172)?
                                    18
                                  :
                                     (X3 <= 224)?
                                      4
                                    :
                                      2
                              :
                                 (X2 <= 171)?
                                  1
                                :
                                  1
              :
                41
            :
               (X1 <= 225)?
                 (X2 <= 213)?
                  2
                :
                   (X1 <= 222)?
                     (X3 <= 224)?
                      3
                    :
                      1
                  :
                    1
              :
                6
    :
       (X1 <= 121)?
        1
      :
         (X3 <= 160)?
          1
        :
           (X1 <= 143)?
            1
          :
             (X1 <= 166)?
              1
            :
              1
;
endmodule
