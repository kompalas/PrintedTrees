module dt(X6, X13, X169, X236, X251, X260, X278, out);
input [-1:0] X6;
input [0:0] X13;
input [1:0] X169;
input [2:0] X236;
input [3:0] X251;
input [4:0] X260;
input [5:0] X278;
output [4:0] out;
assign out = 
   (X278 <= 2)?
    165
  :
     (X278 <= 6)?
      25
    :
       (X278 <= 36)?
         (X13 <= 0)?
          19
        :
           (X278 <= 11)?
            11
          :
             (X169 <= 3)?
              10
            :
               (X6 <= 0)?
                10
              :
                 (X236 <= 4)?
                  4
                :
                   (X251 <= 12)?
                    2
                  :
                    2
      :
         (X278 <= 47)?
          31
        :
           (X260 <= 22)?
            13
          :
            2
;
endmodule
