module top(X0, X1, X2, X3, X4, X5, X6, X7, X8, X9, X10, X11, X12, X13, X14, X15, out);
input [7:0] X0;
input [7:0] X1;
input [7:0] X2;
input [7:0] X3;
input [7:0] X4;
input [7:0] X5;
input [7:0] X6;
input [7:0] X7;
input [7:0] X8;
input [7:0] X9;
input [7:0] X10;
input [7:0] X11;
input [7:0] X12;
input [7:0] X13;
input [7:0] X14;
input [7:0] X15;
output [3:0] out;
assign out = 
   (X15[7:1] <= 34)?
     (X4[7:2] <= 26)?
       (X9[7:1] <= 33)?
         (X14[7:2] <= 35)?
          349
        :
           (X13[7:1] <= 19)?
             (X12 <= 146)?
              19
            :
              21
          :
             (X9[7:3] <= 1)?
              1
            :
              28
      :
         (X5[7:2] <= 46)?
           (X7[7:2] <= 39)?
             (X15[7:1] <= 3)?
               (X5[7:2] <= 8)?
                2
              :
                 (X9[7:1] <= 114)?
                  682
                :
                   (X11[7:2] <= 40)?
                    1
                  :
                    8
            :
               (X5[7:2] <= 40)?
                17
              :
                2
          :
             (X10[7:2] <= 56)?
               (X0[7:3] <= 26)?
                 (X13[7:2] <= 10)?
                   (X12[7:3] <= 22)?
                    1
                  :
                    1
                :
                  21
              :
                 (X13[7:1] <= 49)?
                  4
                :
                  1
            :
              38
        :
           (X9[7:3] <= 21)?
             (X14[7:1] <= 23)?
               (X6[7:2] <= 34)?
                 (X10[7:2] <= 25)?
                   (X7[7:1] <= 72)?
                    1
                  :
                    4
                :
                   (X2[7:2] <= 22)?
                     (X0[7:2] <= 18)?
                      2
                    :
                       (X5 <= 196)?
                        1
                      :
                        1
                  :
                     (X1[7:2] <= 47)?
                      1
                    :
                      91
              :
                 (X9[7:3] <= 16)?
                   (X0[7:2] <= 57)?
                    1
                  :
                    7
                :
                  33
            :
               (X10[7:4] <= 9)?
                 (X12[7:2] <= 34)?
                  19
                :
                   (X7 <= 160)?
                    6
                  :
                    1
              :
                 (X9[7:2] <= 37)?
                   (X13[7:1] <= 17)?
                     (X8[7:4] <= 8)?
                       (X6[7:2] <= 2)?
                        1
                      :
                        1
                    :
                      3
                  :
                    56
                :
                   (X5[7:2] <= 48)?
                    2
                  :
                    7
          :
             (X0[7:2] <= 22)?
               (X7[7:1] <= 115)?
                 (X11[7:2] <= 32)?
                   (X3[7:2] <= 62)?
                    1
                  :
                    3
                :
                  3
              :
                 (X1[7:1] <= 72)?
                  3
                :
                  24
            :
               (X1[7:3] <= 30)?
                207
              :
                 (X7[7:2] <= 38)?
                   (X13 <= 40)?
                    1
                  :
                    5
                :
                   (X5[7:4] <= 16)?
                    29
                  :
                    2
    :
       (X14 <= 146)?
         (X3[7:3] <= 31)?
           (X10[7:3] <= 27)?
             (X7[7:2] <= 34)?
               (X9[7:3] <= 12)?
                13
              :
                 (X5 <= 96)?
                  11
                :
                  1
            :
               (X0[7:2] <= 18)?
                 (X8[7:3] <= 14)?
                   (X13[7:2] <= 19)?
                     (X12[7:1] <= 33)?
                      1
                    :
                       (X1[7:4] <= 9)?
                        1
                      :
                        1
                  :
                    6
                :
                   (X3[7:2] <= 55)?
                     (X2[7:2] <= 6)?
                       (X3[7:1] <= 104)?
                         (X4[7:1] <= 84)?
                          5
                        :
                          1
                      :
                        2
                    :
                       (X13[7:1] <= 61)?
                        211
                      :
                        1
                  :
                     (X2[7:3] <= 13)?
                      9
                    :
                      4
              :
                 (X10[7:3] <= 19)?
                   (X3[7:4] <= 13)?
                     (X5[7:2] <= 44)?
                      2
                    :
                       (X5[7:4] <= 16)?
                        1
                      :
                        1
                  :
                    43
                :
                   (X0[7:4] <= 8)?
                     (X9[7:2] <= 39)?
                      5
                    :
                       (X3[7:2] <= 45)?
                         (X2[7:3] <= 11)?
                          1
                        :
                          1
                      :
                        3
                  :
                     (X7[7:2] <= 46)?
                      1
                    :
                      29
          :
             (X1[7:3] <= 19)?
               (X6[7:4] <= 12)?
                 (X13[7:3] <= 4)?
                  6
                :
                  4
              :
                11
            :
               (X9 <= 83)?
                 (X0[7:3] <= 16)?
                  2
                :
                  3
              :
                 (X0[7:2] <= 4)?
                   (X3[7:3] <= 26)?
                    10
                  :
                     (X2[7:1] <= 60)?
                      3
                    :
                       (X2[7:3] <= 24)?
                        2
                      :
                        1
                :
                   (X9 <= 128)?
                     (X0[7:2] <= 42)?
                      2
                    :
                      5
                  :
                    163
        :
           (X7[7:2] <= 51)?
             (X2[7:2] <= 62)?
               (X4[7:3] <= 17)?
                 (X9[7:3] <= 11)?
                   (X0[7:5] <= 6)?
                    2
                  :
                    7
                :
                   (X6[7:2] <= 49)?
                     (X2[7:2] <= 33)?
                      6
                    :
                       (X14[7:2] <= 20)?
                         (X1[7:1] <= 107)?
                          1
                        :
                           (X10[7:3] <= 10)?
                            1
                          :
                            23
                      :
                        2
                  :
                    9
              :
                 (X12[7:2] <= 17)?
                   (X15[7:1] <= 20)?
                    6
                  :
                     (X13[7:3] <= 1)?
                      1
                    :
                      3
                :
                   (X9[7:1] <= 25)?
                     (X15[7:3] <= 6)?
                      3
                    :
                       (X14[7:3] <= 5)?
                        1
                      :
                        2
                  :
                     (X3[7:1] <= 127)?
                       (X0[7:2] <= 46)?
                         (X6[7:3] <= 32)?
                           (X6[7:4] <= 6)?
                            1
                          :
                            16
                        :
                           (X1 <= 185)?
                            2
                          :
                            3
                      :
                         (X1[7:2] <= 63)?
                          1
                        :
                          3
                    :
                       (X5[7:1] <= 78)?
                        1
                      :
                         (X13[7:2] <= 13)?
                           (X2[7:2] <= 58)?
                            643
                          :
                             (X13[7:4] <= 3)?
                              16
                            :
                              1
                        :
                           (X10[7:4] <= 11)?
                            1
                          :
                            1
            :
               (X5[7:3] <= 27)?
                 (X13[7:3] <= 6)?
                   (X4[7:5] <= 6)?
                     (X2[7:2] <= 61)?
                      2
                    :
                      9
                  :
                     (X10[7:5] <= 3)?
                      2
                    :
                      23
                :
                   (X9[7:3] <= 12)?
                     (X9[7:1] <= 37)?
                      11
                    :
                      1
                  :
                    20
              :
                 (X1[7:1] <= 102)?
                  8
                :
                   (X6[7:3] <= 23)?
                     (X11[7:4] <= 11)?
                      64
                    :
                      1
                  :
                     (X15[7:2] <= 9)?
                       (X11[7:3] <= 9)?
                        1
                      :
                        2
                    :
                      2
          :
             (X5[7:1] <= 115)?
              92
            :
               (X2[7:1] <= 79)?
                 (X11[7:2] <= 27)?
                   (X10[7:2] <= 42)?
                    2
                  :
                    25
                :
                   (X2[7:4] <= 10)?
                    55
                  :
                     (X1[7:2] <= 60)?
                       (X1[7:1] <= 106)?
                        1
                      :
                         (X14[7:1] <= 36)?
                          1
                        :
                          1
                    :
                      4
              :
                 (X13[7:2] <= 11)?
                   (X11[7:3] <= 5)?
                    1
                  :
                    76
                :
                   (X11[7:2] <= 31)?
                    2
                  :
                    1
      :
         (X3[7:2] <= 56)?
           (X6[7:2] <= 21)?
             (X9[7:1] <= 54)?
               (X14[7:5] <= 7)?
                1
              :
                1
            :
              38
          :
             (X8[7:5] <= 3)?
               (X8[7:4] <= 4)?
                6
              :
                1
            :
               (X1[7:2] <= 64)?
                 (X10[7:3] <= 0)?
                   (X6[7:2] <= 58)?
                    12
                  :
                    4
                :
                   (X13[7:2] <= 27)?
                    257
                  :
                    1
              :
                 (X14[7:2] <= 63)?
                  3
                :
                  1
        :
           (X8[7:1] <= 46)?
             (X9[7:1] <= 11)?
               (X8[7:1] <= 18)?
                 (X4[7:1] <= 61)?
                   (X0[7:3] <= 6)?
                    15
                  :
                     (X5[7:1] <= 96)?
                      4
                    :
                      4
                :
                  105
              :
                 (X4[7:3] <= 22)?
                   (X8[7:1] <= 25)?
                     (X7[7:1] <= 39)?
                       (X12[7:2] <= 34)?
                        1
                      :
                        2
                    :
                       (X7[7:2] <= 28)?
                        7
                      :
                        1
                  :
                    15
                :
                   (X1[7:3] <= 28)?
                    26
                  :
                     (X6[7:3] <= 22)?
                      3
                    :
                      1
            :
               (X9[7:2] <= 31)?
                 (X5[7:2] <= 57)?
                  335
                :
                   (X2[7:2] <= 20)?
                    56
                  :
                     (X4[7:4] <= 12)?
                      3
                    :
                      25
              :
                 (X10[7:1] <= 68)?
                  2
                :
                  1
          :
             (X15[7:2] <= 12)?
               (X6 <= 169)?
                 (X2[7:3] <= 10)?
                  18
                :
                   (X13[7:1] <= 11)?
                    80
                  :
                     (X2[7:1] <= 51)?
                      3
                    :
                      7
              :
                 (X8[7:2] <= 48)?
                   (X2[7:3] <= 15)?
                    108
                  :
                     (X4[7:2] <= 55)?
                       (X5[7:1] <= 104)?
                        2
                      :
                        16
                    :
                       (X8[7:2] <= 34)?
                         (X0[7:1] <= 13)?
                           (X2[7:2] <= 34)?
                            2
                          :
                            1
                        :
                          46
                      :
                         (X2[7:3] <= 19)?
                          2
                        :
                          3
                :
                   (X2[7:1] <= 69)?
                     (X14[7:3] <= 24)?
                       (X1[7:3] <= 25)?
                        1
                      :
                        8
                    :
                       (X7[7:2] <= 45)?
                        1
                      :
                        4
                  :
                    15
            :
               (X0[7:3] <= 10)?
                27
              :
                1
  :
     (X13[7:1] <= 76)?
       (X0[7:2] <= 26)?
         (X14[7:3] <= 19)?
           (X1[7:2] <= 54)?
             (X8[7:3] <= 31)?
               (X12[7:2] <= 61)?
                34
              :
                 (X5[7:2] <= 53)?
                  1
                :
                  2
            :
              5
          :
             (X3[7:2] <= 56)?
               (X4 <= 83)?
                2
              :
                8
            :
               (X9[7:2] <= 27)?
                 (X15[7:2] <= 39)?
                  59
                :
                   (X11[7:2] <= 7)?
                    1
                  :
                    1
              :
                2
        :
           (X8[7:2] <= 4)?
             (X0[7:1] <= 14)?
              1
            :
              13
          :
             (X1[7:2] <= 42)?
               (X15[7:4] <= 12)?
                 (X2[7:1] <= 64)?
                  6
                :
                  1
              :
                2
            :
              563
      :
         (X6[7:2] <= 24)?
           (X14[7:4] <= 12)?
             (X9[7:3] <= 11)?
               (X15[7:3] <= 25)?
                324
              :
                1
            :
               (X13[7:1] <= 6)?
                 (X11[7:2] <= 13)?
                  4
                :
                  2
              :
                 (X15[7:1] <= 34)?
                  1
                :
                  12
          :
             (X12 <= 149)?
              17
            :
              29
        :
           (X15[7:1] <= 53)?
             (X7[7:3] <= 15)?
               (X10[7:4] <= 7)?
                 (X2[7:1] <= 42)?
                  1
                :
                  4
              :
                 (X0 <= 134)?
                  2
                :
                  3
            :
               (X11[7:2] <= 10)?
                 (X3 <= 239)?
                   (X4 <= 122)?
                    1
                  :
                    3
                :
                  4
              :
                6
          :
             (X15[7:2] <= 34)?
               (X7[7:2] <= 24)?
                3
              :
                17
            :
              177
    :
       (X8[7:2] <= 38)?
         (X14[7:3] <= 27)?
           (X12[7:2] <= 10)?
            9
          :
             (X11[7:3] <= 10)?
               (X12[7:2] <= 62)?
                16
              :
                12
            :
               (X1[7:3] <= 11)?
                1
              :
                331
        :
           (X13[7:1] <= 96)?
             (X6[7:1] <= 22)?
              4
            :
               (X11[7:1] <= 61)?
                 (X5[7:2] <= 28)?
                   (X9[7:3] <= 5)?
                    1
                  :
                    1
                :
                  40
              :
                 (X5[7:2] <= 43)?
                  3
                :
                  1
          :
             (X12[7:2] <= 55)?
               (X5 <= 143)?
                377
              :
                 (X12[7:4] <= 7)?
                  47
                :
                  1
            :
              1
      :
         (X7 <= 65)?
           (X2[7:2] <= 30)?
             (X6[7:4] <= 16)?
               (X4[7:5] <= 4)?
                716
              :
                 (X3[7:3] <= 17)?
                  1
                :
                  1
            :
               (X15[7:2] <= 54)?
                11
              :
                4
          :
             (X11[7:1] <= 76)?
               (X6[7:2] <= 4)?
                1
              :
                1
            :
              11
        :
           (X9[7:2] <= 41)?
             (X12[7:2] <= 8)?
              1
            :
              31
          :
             (X5[7:2] <= 11)?
               (X6[7:3] <= 17)?
                2
              :
                24
            :
              16
;
endmodule
