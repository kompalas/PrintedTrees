module top(X0, X1, X2, X3, X4, X5, X6, X7, X8, X9, X10, X11, X12, X13, X14, X15, out);
input [7:0] X0;
input [7:0] X1;
input [7:0] X2;
input [7:0] X3;
input [7:0] X4;
input [7:0] X5;
input [7:0] X6;
input [7:0] X7;
input [7:0] X8;
input [7:0] X9;
input [7:0] X10;
input [7:0] X11;
input [7:0] X12;
input [7:0] X13;
input [7:0] X14;
input [7:0] X15;
output [3:0] out;
assign out = 
   (X15 <= 63)?
     (X4 <= 104)?
       (X9 <= 55)?
         (X14 <= 133)?
          349
        :
           (X13 <= 38)?
             (X12 <= 143)?
              19
            :
              21
          :
             (X9 <= 19)?
              1
            :
              28
      :
         (X5 <= 170)?
           (X7 <= 155)?
             (X15 <= 3)?
               (X5 <= 23)?
                2
              :
                 (X9 <= 227)?
                  682
                :
                   (X11 <= 159)?
                    1
                  :
                    8
            :
               (X5 <= 143)?
                17
              :
                2
          :
             (X10 <= 210)?
               (X0 <= 196)?
                 (X13 <= 28)?
                   (X12 <= 148)?
                    1
                  :
                    1
                :
                  21
              :
                 (X13 <= 93)?
                  4
                :
                  1
            :
              38
        :
           (X9 <= 160)?
             (X14 <= 42)?
               (X6 <= 127)?
                 (X10 <= 88)?
                   (X7 <= 140)?
                    1
                  :
                    4
                :
                   (X2 <= 79)?
                     (X0 <= 69)?
                      2
                    :
                       (X5 <= 193)?
                        1
                      :
                        1
                  :
                     (X1 <= 195)?
                      1
                    :
                      91
              :
                 (X9 <= 120)?
                   (X0 <= 221)?
                    1
                  :
                    7
                :
                  33
            :
               (X10 <= 111)?
                 (X12 <= 131)?
                  19
                :
                   (X7 <= 156)?
                    6
                  :
                    1
              :
                 (X9 <= 143)?
                   (X13 <= 37)?
                     (X8 <= 124)?
                       (X6 <= 9)?
                        1
                      :
                        1
                    :
                      3
                  :
                    56
                :
                   (X5 <= 183)?
                    2
                  :
                    7
          :
             (X0 <= 83)?
               (X7 <= 228)?
                 (X11 <= 118)?
                   (X3 <= 243)?
                    1
                  :
                    3
                :
                  3
              :
                 (X1 <= 138)?
                  3
                :
                  24
            :
               (X1 <= 237)?
                207
              :
                 (X7 <= 160)?
                   (X13 <= 38)?
                    1
                  :
                    5
                :
                   (X5 <= 227)?
                    29
                  :
                    2
    :
       (X14 <= 145)?
         (X3 <= 234)?
           (X10 <= 209)?
             (X7 <= 137)?
               (X9 <= 81)?
                13
              :
                 (X5 <= 97)?
                  11
                :
                  1
            :
               (X0 <= 51)?
                 (X8 <= 101)?
                   (X13 <= 58)?
                     (X12 <= 67)?
                      1
                    :
                       (X1 <= 111)?
                        1
                      :
                        1
                  :
                    6
                :
                   (X3 <= 219)?
                     (X2 <= 6)?
                       (X3 <= 198)?
                         (X4 <= 157)?
                          5
                        :
                          1
                      :
                        2
                    :
                       (X13 <= 116)?
                        211
                      :
                        1
                  :
                     (X2 <= 84)?
                      9
                    :
                      4
              :
                 (X10 <= 148)?
                   (X3 <= 196)?
                     (X5 <= 174)?
                      2
                    :
                       (X5 <= 219)?
                        1
                      :
                        1
                  :
                    43
                :
                   (X0 <= 90)?
                     (X9 <= 150)?
                      5
                    :
                       (X3 <= 170)?
                         (X2 <= 82)?
                          1
                        :
                          1
                      :
                        3
                  :
                     (X7 <= 174)?
                      1
                    :
                      29
          :
             (X1 <= 142)?
               (X6 <= 133)?
                 (X13 <= 35)?
                  6
                :
                  4
              :
                11
            :
               (X9 <= 81)?
                 (X0 <= 124)?
                  2
                :
                  3
              :
                 (X0 <= 3)?
                   (X3 <= 195)?
                    10
                  :
                     (X2 <= 124)?
                      3
                    :
                       (X2 <= 173)?
                        2
                      :
                        1
                :
                   (X9 <= 124)?
                     (X0 <= 180)?
                      2
                    :
                      5
                  :
                    163
        :
           (X7 <= 196)?
             (X2 <= 229)?
               (X4 <= 137)?
                 (X9 <= 67)?
                   (X0 <= 128)?
                    2
                  :
                    7
                :
                   (X6 <= 183)?
                     (X2 <= 123)?
                      6
                    :
                       (X14 <= 64)?
                         (X1 <= 212)?
                          1
                        :
                           (X10 <= 68)?
                            1
                          :
                            23
                      :
                        2
                  :
                    9
              :
                 (X12 <= 64)?
                   (X15 <= 36)?
                    6
                  :
                     (X13 <= 4)?
                      1
                    :
                      3
                :
                   (X9 <= 47)?
                     (X15 <= 42)?
                      3
                    :
                       (X14 <= 40)?
                        1
                      :
                        2
                  :
                     (X3 <= 250)?
                       (X0 <= 182)?
                         (X6 <= 225)?
                           (X6 <= 96)?
                            1
                          :
                            16
                        :
                           (X1 <= 182)?
                            2
                          :
                            3
                      :
                         (X1 <= 248)?
                          1
                        :
                          3
                    :
                       (X5 <= 156)?
                        1
                      :
                         (X13 <= 42)?
                           (X2 <= 221)?
                            643
                          :
                             (X13 <= 9)?
                              16
                            :
                              1
                        :
                           (X10 <= 180)?
                            1
                          :
                            1
            :
               (X5 <= 219)?
                 (X13 <= 27)?
                   (X4 <= 197)?
                     (X2 <= 243)?
                      2
                    :
                      9
                  :
                     (X10 <= 95)?
                      2
                    :
                      23
                :
                   (X9 <= 99)?
                     (X9 <= 67)?
                      11
                    :
                      1
                  :
                    20
              :
                 (X1 <= 205)?
                  8
                :
                   (X6 <= 152)?
                     (X11 <= 127)?
                      64
                    :
                      1
                  :
                     (X15 <= 19)?
                       (X11 <= 73)?
                        1
                      :
                        2
                    :
                      2
          :
             (X5 <= 229)?
              92
            :
               (X2 <= 150)?
                 (X11 <= 97)?
                   (X10 <= 152)?
                    2
                  :
                    25
                :
                   (X2 <= 104)?
                    55
                  :
                     (X1 <= 241)?
                       (X1 <= 212)?
                        1
                      :
                         (X14 <= 74)?
                          1
                        :
                          1
                    :
                      4
              :
                 (X13 <= 46)?
                   (X11 <= 38)?
                    1
                  :
                    76
                :
                   (X11 <= 123)?
                    2
                  :
                    1
      :
         (X3 <= 224)?
           (X6 <= 84)?
             (X9 <= 109)?
               (X14 <= 253)?
                1
              :
                1
            :
              38
          :
             (X8 <= 68)?
               (X8 <= 64)?
                6
              :
                1
            :
               (X1 <= 238)?
                 (X10 <= 1)?
                   (X6 <= 214)?
                    12
                  :
                    4
                :
                   (X13 <= 104)?
                    257
                  :
                    1
              :
                 (X14 <= 239)?
                  3
                :
                  1
        :
           (X8 <= 88)?
             (X9 <= 22)?
               (X8 <= 32)?
                 (X4 <= 122)?
                   (X0 <= 32)?
                    15
                  :
                     (X5 <= 183)?
                      4
                    :
                      4
                :
                  105
              :
                 (X4 <= 168)?
                   (X8 <= 50)?
                     (X7 <= 74)?
                       (X12 <= 127)?
                        1
                      :
                        2
                    :
                       (X7 <= 116)?
                        7
                      :
                        1
                  :
                    15
                :
                   (X1 <= 230)?
                    26
                  :
                     (X6 <= 160)?
                      3
                    :
                      1
            :
               (X9 <= 124)?
                 (X5 <= 224)?
                  335
                :
                   (X2 <= 81)?
                    56
                  :
                     (X4 <= 155)?
                      3
                    :
                      25
              :
                 (X10 <= 137)?
                  2
                :
                  1
          :
             (X15 <= 40)?
               (X6 <= 165)?
                 (X2 <= 73)?
                  18
                :
                   (X13 <= 20)?
                    80
                  :
                     (X2 <= 105)?
                      3
                    :
                      7
              :
                 (X8 <= 183)?
                   (X2 <= 124)?
                    108
                  :
                     (X4 <= 221)?
                       (X5 <= 202)?
                        2
                      :
                        16
                    :
                       (X8 <= 134)?
                         (X0 <= 19)?
                           (X2 <= 137)?
                            2
                          :
                            1
                        :
                          46
                      :
                         (X2 <= 140)?
                          2
                        :
                          3
                :
                   (X2 <= 136)?
                     (X14 <= 189)?
                       (X1 <= 174)?
                        1
                      :
                        8
                    :
                       (X7 <= 182)?
                        1
                      :
                        4
                  :
                    15
            :
               (X0 <= 73)?
                27
              :
                1
  :
     (X13 <= 152)?
       (X0 <= 91)?
         (X14 <= 127)?
           (X1 <= 216)?
             (X8 <= 223)?
               (X12 <= 237)?
                34
              :
                 (X5 <= 210)?
                  1
                :
                  2
            :
              5
          :
             (X3 <= 215)?
               (X4 <= 81)?
                2
              :
                8
            :
               (X9 <= 92)?
                 (X15 <= 151)?
                  59
                :
                   (X11 <= 27)?
                    1
                  :
                    1
              :
                2
        :
           (X8 <= 3)?
             (X0 <= 19)?
              1
            :
              13
          :
             (X1 <= 178)?
               (X15 <= 165)?
                 (X2 <= 124)?
                  6
                :
                  1
              :
                2
            :
              563
      :
         (X6 <= 78)?
           (X14 <= 168)?
             (X9 <= 76)?
               (X15 <= 200)?
                324
              :
                1
            :
               (X13 <= 13)?
                 (X11 <= 51)?
                  4
                :
                  2
              :
                 (X15 <= 65)?
                  1
                :
                  12
          :
             (X12 <= 147)?
              17
            :
              29
        :
           (X15 <= 104)?
             (X7 <= 116)?
               (X10 <= 82)?
                 (X2 <= 83)?
                  1
                :
                  4
              :
                 (X0 <= 132)?
                  2
                :
                  3
            :
               (X11 <= 22)?
                 (X3 <= 239)?
                   (X4 <= 120)?
                    1
                  :
                    3
                :
                  4
              :
                6
          :
             (X15 <= 134)?
               (X7 <= 87)?
                3
              :
                17
            :
              177
    :
       (X8 <= 134)?
         (X14 <= 214)?
           (X12 <= 40)?
            9
          :
             (X11 <= 81)?
               (X12 <= 238)?
                16
              :
                12
            :
               (X1 <= 90)?
                1
              :
                331
        :
           (X13 <= 191)?
             (X6 <= 36)?
              4
            :
               (X11 <= 116)?
                 (X5 <= 97)?
                   (X9 <= 10)?
                    1
                  :
                    1
                :
                  40
              :
                 (X5 <= 165)?
                  3
                :
                  1
          :
             (X12 <= 211)?
               (X5 <= 140)?
                377
              :
                 (X12 <= 111)?
                  47
                :
                  1
            :
              1
      :
         (X7 <= 63)?
           (X2 <= 129)?
             (X6 <= 250)?
               (X4 <= 142)?
                716
              :
                 (X3 <= 118)?
                  1
                :
                  1
            :
               (X15 <= 216)?
                11
              :
                4
          :
             (X11 <= 142)?
               (X6 <= 13)?
                1
              :
                1
            :
              11
        :
           (X9 <= 150)?
             (X12 <= 32)?
              1
            :
              31
          :
             (X5 <= 42)?
               (X6 <= 124)?
                2
              :
                24
            :
              16
;
endmodule
