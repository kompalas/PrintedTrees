module top(X0, X1, X2, X3, X4, X5, X6, X7, X8, X9, X10, out);
input [7:0] X0;
input [7:0] X1;
input [7:0] X2;
input [7:0] X3;
input [7:0] X4;
input [7:0] X5;
input [7:0] X6;
input [7:0] X7;
input [7:0] X8;
input [7:0] X9;
input [7:0] X10;
output [3:0] out;
assign out = 
   (X10[7:3] <= 9)?
     (X0[7:2] <= 37)?
       (X6[7:2] <= 22)?
         (X9[7:1] <= 17)?
           (X3[7:3] <= 11)?
             (X4[7:1] <= 12)?
               (X6[7:2] <= 19)?
                 (X2[7:1] <= 41)?
                   (X9[7:1] <= 15)?
                     (X0[7:2] <= 21)?
                       (X9[7:4] <= 4)?
                        13
                      :
                         (X0[7:5] <= 2)?
                           (X4[7:2] <= 10)?
                            1
                          :
                            5
                        :
                          2
                    :
                       (X10[7:1] <= 29)?
                        1
                      :
                        2
                  :
                    20
                :
                   (X1[7:3] <= 3)?
                    1
                  :
                     (X9[7:2] <= 7)?
                      1
                    :
                      4
              :
                3
            :
               (X4[7:3] <= 10)?
                 (X7[7:1] <= 70)?
                  20
                :
                   (X7[7:3] <= 18)?
                     (X0[7:2] <= 19)?
                      2
                    :
                      3
                  :
                    12
              :
                1
          :
             (X2[7:1] <= 17)?
              1
            :
              3
        :
           (X1[7:1] <= 48)?
             (X1[7:2] <= 6)?
              5
            :
               (X0[7:2] <= 24)?
                 (X1[7:2] <= 12)?
                   (X7[7:1] <= 59)?
                    3
                  :
                     (X6[7:3] <= 10)?
                       (X1[7:3] <= 11)?
                        7
                      :
                         (X10[7:4] <= 4)?
                          1
                        :
                          1
                    :
                      1
                :
                   (X0 <= 45)?
                    11
                  :
                     (X2[7:3] <= 1)?
                      8
                    :
                       (X6 <= 31)?
                         (X7[7:3] <= 14)?
                          7
                        :
                           (X7[7:2] <= 36)?
                             (X0[7:5] <= 2)?
                               (X4[7:3] <= 8)?
                                 (X8[7:2] <= 29)?
                                  11
                                :
                                   (X8[7:2] <= 34)?
                                    3
                                  :
                                     (X10[7:5] <= 1)?
                                      1
                                    :
                                       (X9[7:2] <= 16)?
                                        1
                                      :
                                        7
                              :
                                2
                            :
                              3
                          :
                             (X8[7:3] <= 14)?
                               (X7[7:2] <= 36)?
                                1
                              :
                                1
                            :
                              8
                      :
                         (X3[7:5] <= 0)?
                          14
                        :
                           (X0[7:2] <= 18)?
                             (X4[7:2] <= 8)?
                               (X4[7:1] <= 17)?
                                 (X1[7:1] <= 24)?
                                  1
                                :
                                  13
                              :
                                 (X1[7:1] <= 42)?
                                   (X2[7:4] <= 9)?
                                     (X1[7:1] <= 33)?
                                      2
                                    :
                                       (X0[7:2] <= 18)?
                                        3
                                      :
                                        1
                                  :
                                    4
                                :
                                  7
                            :
                              10
                          :
                             (X9[7:4] <= 2)?
                              1
                            :
                              8
              :
                 (X0[7:2] <= 31)?
                   (X9[7:2] <= 11)?
                     (X9[7:2] <= 14)?
                      18
                    :
                       (X0[7:2] <= 32)?
                        1
                      :
                        1
                  :
                     (X0[7:2] <= 26)?
                       (X9 <= 51)?
                        3
                      :
                         (X9[7:3] <= 20)?
                          7
                        :
                          1
                    :
                       (X7[7:3] <= 30)?
                        13
                      :
                         (X1[7:2] <= 16)?
                          1
                        :
                          2
                :
                   (X2[7:2] <= 34)?
                     (X0[7:1] <= 66)?
                      7
                    :
                      1
                  :
                    5
          :
             (X10[7:2] <= 10)?
              2
            :
               (X1[7:4] <= 10)?
                 (X0 <= 101)?
                   (X8[7:2] <= 28)?
                     (X5[7:3] <= 6)?
                       (X10[7:3] <= 7)?
                        2
                      :
                        1
                    :
                      8
                  :
                     (X7[7:3] <= 15)?
                       (X9[7:2] <= 8)?
                         (X5[7:2] <= 8)?
                          2
                        :
                          3
                      :
                         (X0[7:2] <= 11)?
                           (X4[7:5] <= 0)?
                             (X7[7:3] <= 17)?
                              6
                            :
                              1
                          :
                            2
                        :
                          13
                    :
                      13
                :
                   (X10 <= 46)?
                    3
                  :
                     (X2[7:1] <= 16)?
                      1
                    :
                      1
              :
                 (X9[7:3] <= 10)?
                  2
                :
                  2
      :
         (X4[7:4] <= 1)?
           (X6[7:4] <= 6)?
            2
          :
            3
        :
          45
    :
       (X9[7:1] <= 23)?
         (X1[7:2] <= 18)?
          5
        :
          1
      :
         (X5[7:3] <= 9)?
           (X9[7:3] <= 11)?
            13
          :
             (X0[7:4] <= 15)?
               (X9[7:3] <= 11)?
                1
              :
                3
            :
               (X7[7:2] <= 45)?
                1
              :
                2
        :
          2
  :
     (X9[7:3] <= 8)?
       (X10[7:2] <= 33)?
         (X6[7:2] <= 6)?
           (X1[7:4] <= 7)?
             (X3[7:2] <= 3)?
               (X8[7:4] <= 10)?
                 (X7[7:1] <= 59)?
                  5
                :
                   (X8[7:3] <= 14)?
                    1
                  :
                    2
              :
                 (X2[7:4] <= 0)?
                   (X8[7:5] <= 4)?
                    2
                  :
                     (X3[7:3] <= 3)?
                      1
                    :
                      1
                :
                  7
            :
               (X9 <= 39)?
                 (X1[7:4] <= 5)?
                   (X3[7:1] <= 14)?
                    5
                  :
                     (X0[7:3] <= 9)?
                       (X9[7:3] <= 4)?
                        4
                      :
                        2
                    :
                       (X0[7:1] <= 41)?
                        4
                      :
                         (X8[7:2] <= 27)?
                          6
                        :
                          1
                :
                   (X4[7:4] <= 5)?
                     (X6[7:3] <= 0)?
                      1
                    :
                       (X5[7:5] <= 2)?
                        15
                      :
                        1
                  :
                    1
              :
                 (X4[7:1] <= 15)?
                   (X10 <= 89)?
                    4
                  :
                     (X0[7:3] <= 16)?
                      1
                    :
                      1
                :
                   (X0[7:3] <= 20)?
                     (X6[7:1] <= 10)?
                      9
                    :
                      1
                  :
                    1
          :
             (X9[7:1] <= 14)?
               (X6[7:4] <= 3)?
                 (X1[7:4] <= 15)?
                   (X1[7:3] <= 17)?
                    1
                  :
                    3
                :
                  2
              :
                1
            :
               (X2[7:3] <= 4)?
                3
              :
                 (X7[7:2] <= 32)?
                  3
                :
                  1
        :
           (X9[7:3] <= 4)?
             (X10[7:1] <= 55)?
               (X3[7:2] <= 11)?
                 (X3[7:2] <= 6)?
                   (X4[7:4] <= 4)?
                    4
                  :
                    8
                :
                  25
              :
                 (X10[7:3] <= 13)?
                  2
                :
                  4
            :
               (X5[7:2] <= 21)?
                 (X2[7:2] <= 5)?
                   (X2[7:2] <= 0)?
                    1
                  :
                    2
                :
                  2
              :
                1
          :
             (X7[7:1] <= 75)?
               (X0[7:2] <= 25)?
                 (X1[7:1] <= 25)?
                   (X10[7:2] <= 17)?
                    1
                  :
                    4
                :
                   (X2[7:3] <= 3)?
                     (X5[7:1] <= 63)?
                       (X0 <= 78)?
                        19
                      :
                        1
                    :
                      2
                  :
                     (X2[7:3] <= 12)?
                       (X9 <= 43)?
                        8
                      :
                         (X6[7:2] <= 13)?
                          1
                        :
                          2
                    :
                       (X9[7:3] <= 6)?
                         (X5[7:4] <= 6)?
                           (X3[7:1] <= 13)?
                            4
                          :
                            3
                        :
                          9
                      :
                        2
              :
                 (X0[7:3] <= 12)?
                  1
                :
                  6
            :
              10
      :
         (X1[7:3] <= 8)?
           (X3[7:4] <= 5)?
             (X2[7:2] <= 43)?
               (X0[7:2] <= 2)?
                1
              :
                 (X4 <= 7)?
                  2
                :
                   (X6[7:3] <= 4)?
                     (X0[7:2] <= 29)?
                       (X0[7:4] <= 4)?
                         (X6[7:2] <= 4)?
                          1
                        :
                           (X6[7:5] <= 1)?
                            9
                          :
                             (X7[7:3] <= 11)?
                              1
                            :
                              1
                      :
                        3
                    :
                      8
                  :
                    20
            :
               (X8[7:2] <= 26)?
                1
              :
                1
          :
             (X2[7:3] <= 14)?
               (X7[7:5] <= 3)?
                1
              :
                2
            :
              5
        :
           (X7 <= 70)?
             (X8 <= 215)?
               (X2[7:3] <= 2)?
                 (X9[7:3] <= 8)?
                  3
                :
                  2
              :
                6
            :
              2
          :
             (X1[7:3] <= 14)?
               (X1 <= 85)?
                1
              :
                 (X4[7:3] <= 1)?
                  1
                :
                  7
            :
               (X1[7:5] <= 5)?
                1
              :
                1
    :
       (X10[7:1] <= 61)?
         (X1[7:2] <= 11)?
           (X6[7:4] <= 6)?
             (X8[7:2] <= 26)?
               (X0[7:1] <= 35)?
                 (X7[7:3] <= 14)?
                   (X10[7:2] <= 32)?
                    1
                  :
                    1
                :
                  2
              :
                 (X2[7:3] <= 21)?
                   (X3[7:2] <= 11)?
                     (X3[7:3] <= 6)?
                       (X6[7:3] <= 4)?
                         (X10[7:2] <= 22)?
                          7
                        :
                           (X1[7:2] <= 7)?
                            1
                          :
                            3
                      :
                         (X0[7:1] <= 53)?
                          3
                        :
                           (X7 <= 164)?
                             (X7[7:4] <= 7)?
                               (X2[7:2] <= 29)?
                                3
                              :
                                2
                            :
                              11
                          :
                            1
                    :
                       (X8[7:3] <= 9)?
                        1
                      :
                        1
                  :
                    6
                :
                  5
            :
               (X5[7:3] <= 5)?
                 (X9[7:2] <= 19)?
                   (X2 <= 94)?
                    3
                  :
                     (X2[7:4] <= 11)?
                       (X6[7:2] <= 2)?
                        1
                      :
                         (X6[7:3] <= 1)?
                           (X4[7:4] <= 2)?
                            2
                          :
                            1
                        :
                          2
                    :
                      5
                :
                   (X2[7:2] <= 37)?
                    8
                  :
                    1
              :
                 (X9[7:4] <= 9)?
                  10
                :
                   (X7[7:2] <= 28)?
                    5
                  :
                     (X7[7:4] <= 10)?
                       (X1[7:4] <= 4)?
                         (X10[7:2] <= 21)?
                          2
                        :
                          2
                      :
                        6
                    :
                      2
          :
             (X5[7:2] <= 31)?
               (X2[7:1] <= 73)?
                 (X8[7:4] <= 10)?
                  8
                :
                   (X2[7:3] <= 16)?
                    5
                  :
                    2
              :
                3
            :
               (X0[7:3] <= 10)?
                4
              :
                5
        :
           (X6 <= 66)?
             (X4[7:4] <= 4)?
               (X1[7:2] <= 26)?
                 (X1[7:3] <= 7)?
                   (X7[7:1] <= 68)?
                     (X7[7:4] <= 10)?
                       (X9[7:2] <= 18)?
                        8
                      :
                         (X7[7:5] <= 1)?
                          2
                        :
                          1
                    :
                      2
                  :
                     (X9[7:3] <= 8)?
                      1
                    :
                      12
                :
                   (X0[7:4] <= 3)?
                     (X8[7:3] <= 25)?
                      17
                    :
                      1
                  :
                     (X1 <= 65)?
                      3
                    :
                       (X8[7:3] <= 9)?
                        3
                      :
                         (X8[7:4] <= 12)?
                          20
                        :
                           (X2[7:3] <= 1)?
                            6
                          :
                            6
              :
                 (X1[7:4] <= 5)?
                  4
                :
                   (X10 <= 81)?
                     (X7[7:2] <= 38)?
                      5
                    :
                      3
                  :
                     (X1 <= 138)?
                      11
                    :
                      1
            :
               (X6[7:3] <= 6)?
                 (X2[7:2] <= 15)?
                   (X3 <= 26)?
                    2
                  :
                     (X3 <= 51)?
                       (X3[7:3] <= 4)?
                        4
                      :
                         (X5[7:2] <= 23)?
                          1
                        :
                          1
                    :
                      1
                :
                   (X2[7:5] <= 5)?
                     (X4[7:3] <= 8)?
                      12
                    :
                      1
                  :
                    2
              :
                6
          :
             (X9 <= 132)?
               (X2[7:2] <= 15)?
                 (X3[7:1] <= 11)?
                  1
                :
                   (X10[7:4] <= 10)?
                    1
                  :
                    1
              :
                15
            :
              4
      :
         (X10[7:4] <= 13)?
           (X9 <= 57)?
             (X6 <= 10)?
               (X3[7:3] <= 6)?
                1
              :
                6
            :
               (X3[7:3] <= 6)?
                 (X2[7:3] <= 16)?
                  1
                :
                  1
              :
                 (X0 <= 181)?
                   (X9[7:6] <= 4)?
                    14
                  :
                    1
                :
                  1
          :
             (X5[7:4] <= 6)?
               (X9[7:2] <= 20)?
                 (X0 <= 127)?
                  22
                :
                   (X3[7:3] <= 4)?
                    1
                  :
                    3
              :
                 (X5[7:2] <= 7)?
                   (X1[7:3] <= 9)?
                    1
                  :
                    5
                :
                  3
            :
               (X3[7:2] <= 11)?
                 (X10[7:3] <= 16)?
                  4
                :
                   (X2 <= 14)?
                    3
                  :
                     (X6[7:1] <= 14)?
                      4
                    :
                       (X6[7:1] <= 18)?
                        3
                      :
                         (X4[7:5] <= 0)?
                          2
                        :
                           (X8[7:3] <= 15)?
                             (X10[7:3] <= 20)?
                              2
                            :
                               (X4[7:1] <= 17)?
                                2
                              :
                                1
                          :
                            6
              :
                 (X10[7:1] <= 87)?
                  3
                :
                  1
        :
           (X6[7:4] <= 2)?
             (X4[7:2] <= 6)?
              2
            :
               (X9 <= 67)?
                3
              :
                2
          :
             (X5[7:5] <= 2)?
              2
            :
              3
;
endmodule
