module top(X0, X1, X4, X5, X6, out);
input [7:0] X0;
input [7:0] X1;
input [7:0] X4;
input [7:0] X5;
input [7:0] X6;
output [1:0] out;
assign out = 
   (X6[7:6] <= 2)?
     (X0[7:4] <= 5)?
       (X6[7:6] <= 1)?
         (X5[7:5] <= 3)?
          3
        :
           (X1[7:6] <= 2)?
            6
          :
            1
      :
        43
    :
       (X5[7:6] <= 4)?
         (X4[7:5] <= 7)?
          37
        :
           (X5[7:6] <= 1)?
            5
          :
            2
      :
        2
  :
     (X5[7:6] <= 1)?
       (X1[7:6] <= 2)?
        1
      :
        3
    :
      44
;
endmodule
