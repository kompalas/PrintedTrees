module top(X0, X1, X4, X5, X6, out);
input [7:0] X0;
input [7:0] X1;
input [7:0] X4;
input [7:0] X5;
input [7:0] X6;
output [1:0] out;
assign out = 
   (X6[7:3] <= 15)?
     (X0[7:4] <= 5)?
       (X6[7:3] <= 9)?
         (X5[7:4] <= 7)?
          3
        :
           (X1[7:5] <= 3)?
            6
          :
            1
      :
        43
    :
       (X5[7:5] <= 7)?
         (X4[7:6] <= 4)?
          37
        :
           (X5[7:4] <= 7)?
            5
          :
            2
      :
        2
  :
     (X5[7:6] <= 1)?
       (X1[7:5] <= 6)?
        1
      :
        3
    :
      44
;
endmodule
