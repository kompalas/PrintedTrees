module top(X561, out);
input [7:0] X561;
output [2:0] out;
assign out = 
   (X561[7:4] <= 7)?
    542
  :
     (X561[7:4] <= 11)?
       (X561[7:4] <= 7)?
         (X561[7:4] <= 7)?
          455
        :
          477
      :
        575
    :
       (X561[7:4] <= 11)?
        545
      :
        382
;
endmodule
