module top(X0, X1, X2, X3, X4, X5, out);
input [7:0] X0;
input [7:0] X1;
input [7:0] X2;
input [7:0] X3;
input [7:0] X4;
input [7:0] X5;
output [1:0] out;
assign out = 
   (X5 <= 17)?
     (X3 <= 52)?
       (X4 <= 128)?
        13
      :
         (X1 <= 79)?
           (X0 <= 16)?
            1
          :
            11
        :
           (X4 <= 153)?
             (X1 <= 130)?
               (X0 <= 48)?
                 (X5 <= 10)?
                  8
                :
                   (X4 <= 151)?
                    1
                  :
                    1
              :
                 (X3 <= 47)?
                  3
                :
                   (X0 <= 54)?
                    1
                  :
                    4
            :
              6
          :
             (X5 <= 8)?
               (X1 <= 114)?
                7
              :
                1
            :
              2
    :
       (X4 <= 128)?
         (X3 <= 80)?
           (X1 <= 147)?
             (X4 <= 112)?
              6
            :
               (X5 <= 8)?
                 (X5 <= 3)?
                  1
                :
                  3
              :
                3
          :
             (X2 <= 85)?
              1
            :
              2
        :
           (X0 <= 115)?
             (X0 <= 110)?
              2
            :
              2
          :
            5
      :
        29
  :
     (X5 <= 25)?
       (X5 <= 25)?
         (X4 <= 142)?
          24
        :
           (X2 <= 86)?
            3
          :
            1
      :
        1
    :
      75
;
endmodule
