module top(X0, X1, X2, X3, X4, X5, X6, X7, X8, X9, X10, out);
input [7:0] X0;
input [7:0] X1;
input [7:0] X2;
input [7:0] X3;
input [7:0] X4;
input [7:0] X5;
input [7:0] X6;
input [7:0] X7;
input [7:0] X8;
input [7:0] X9;
input [7:0] X10;
output [3:0] out;
assign out = 
   (X10 <= 57)?
     (X0 <= 139)?
       (X6 <= 84)?
         (X9 <= 31)?
           (X3 <= 60)?
             (X4 <= 30)?
               (X6 <= 75)?
                 (X2 <= 79)?
                   (X9 <= 24)?
                     (X0 <= 84)?
                       (X9 <= 22)?
                        13
                      :
                         (X0 <= 60)?
                           (X4 <= 25)?
                            1
                          :
                            5
                        :
                          2
                    :
                       (X10 <= 49)?
                        1
                      :
                        2
                  :
                    20
                :
                   (X1 <= 26)?
                    1
                  :
                     (X9 <= 21)?
                      1
                    :
                      4
              :
                3
            :
               (X4 <= 76)?
                 (X7 <= 139)?
                  20
                :
                   (X7 <= 145)?
                     (X0 <= 76)?
                      2
                    :
                      3
                  :
                    12
              :
                1
          :
             (X2 <= 26)?
              1
            :
              3
        :
           (X1 <= 92)?
             (X1 <= 29)?
              5
            :
               (X0 <= 89)?
                 (X1 <= 46)?
                   (X7 <= 118)?
                    3
                  :
                     (X6 <= 64)?
                       (X1 <= 45)?
                        7
                      :
                         (X10 <= 47)?
                          1
                        :
                          1
                    :
                      1
                :
                   (X0 <= 44)?
                    11
                  :
                     (X2 <= 1)?
                      8
                    :
                       (X6 <= 29)?
                         (X7 <= 110)?
                          7
                        :
                           (X7 <= 141)?
                             (X0 <= 76)?
                               (X4 <= 68)?
                                 (X8 <= 115)?
                                  11
                                :
                                   (X8 <= 125)?
                                    3
                                  :
                                     (X10 <= 41)?
                                      1
                                    :
                                       (X9 <= 46)?
                                        1
                                      :
                                        7
                              :
                                2
                            :
                              3
                          :
                             (X8 <= 110)?
                               (X7 <= 151)?
                                1
                              :
                                1
                            :
                              8
                      :
                         (X3 <= 15)?
                          14
                        :
                           (X0 <= 74)?
                             (X4 <= 34)?
                               (X4 <= 28)?
                                 (X1 <= 51)?
                                  1
                                :
                                  13
                              :
                                 (X1 <= 83)?
                                   (X2 <= 83)?
                                     (X1 <= 60)?
                                      2
                                    :
                                       (X0 <= 71)?
                                        3
                                      :
                                        1
                                  :
                                    4
                                :
                                  7
                            :
                              10
                          :
                             (X9 <= 35)?
                              1
                            :
                              8
              :
                 (X0 <= 123)?
                   (X9 <= 42)?
                     (X9 <= 41)?
                      18
                    :
                       (X0 <= 110)?
                        1
                      :
                        1
                  :
                     (X0 <= 101)?
                       (X9 <= 47)?
                        3
                      :
                         (X9 <= 162)?
                          7
                        :
                          1
                    :
                       (X7 <= 206)?
                        13
                      :
                         (X1 <= 66)?
                          1
                        :
                          2
                :
                   (X2 <= 128)?
                     (X0 <= 134)?
                      7
                    :
                      1
                  :
                    5
          :
             (X10 <= 26)?
              2
            :
               (X1 <= 129)?
                 (X0 <= 101)?
                   (X8 <= 94)?
                     (X5 <= 38)?
                       (X10 <= 35)?
                        2
                      :
                        1
                    :
                      8
                  :
                     (X7 <= 135)?
                       (X9 <= 33)?
                         (X5 <= 32)?
                          2
                        :
                          3
                      :
                         (X0 <= 56)?
                           (X4 <= 40)?
                             (X7 <= 132)?
                              6
                            :
                              1
                          :
                            2
                        :
                          13
                    :
                      13
                :
                   (X10 <= 45)?
                    3
                  :
                     (X2 <= 24)?
                      1
                    :
                      1
              :
                 (X9 <= 38)?
                  2
                :
                  2
      :
         (X4 <= 26)?
           (X6 <= 100)?
            2
          :
            3
        :
          45
    :
       (X9 <= 38)?
         (X1 <= 74)?
          5
        :
          1
      :
         (X5 <= 61)?
           (X9 <= 71)?
            13
          :
             (X0 <= 176)?
               (X9 <= 74)?
                1
              :
                3
            :
               (X7 <= 172)?
                1
              :
                2
        :
          2
  :
     (X9 <= 45)?
       (X10 <= 120)?
         (X6 <= 21)?
           (X1 <= 116)?
             (X3 <= 17)?
               (X8 <= 120)?
                 (X7 <= 118)?
                  5
                :
                   (X8 <= 77)?
                    1
                  :
                    2
              :
                 (X2 <= 9)?
                   (X8 <= 133)?
                    2
                  :
                     (X3 <= 12)?
                      1
                    :
                      1
                :
                  7
            :
               (X9 <= 39)?
                 (X1 <= 82)?
                   (X3 <= 20)?
                    5
                  :
                     (X0 <= 63)?
                       (X9 <= 34)?
                        4
                      :
                        2
                    :
                       (X0 <= 86)?
                        4
                      :
                         (X8 <= 109)?
                          6
                        :
                          1
                :
                   (X4 <= 43)?
                     (X6 <= 4)?
                      1
                    :
                       (X5 <= 49)?
                        15
                      :
                        1
                  :
                    1
              :
                 (X4 <= 29)?
                   (X10 <= 87)?
                    4
                  :
                     (X0 <= 106)?
                      1
                    :
                      1
                :
                   (X0 <= 127)?
                     (X6 <= 19)?
                      9
                    :
                      1
                  :
                    1
          :
             (X9 <= 31)?
               (X6 <= 12)?
                 (X1 <= 156)?
                   (X1 <= 133)?
                    1
                  :
                    3
                :
                  2
              :
                1
            :
               (X2 <= 4)?
                3
              :
                 (X7 <= 117)?
                  3
                :
                  1
        :
           (X9 <= 31)?
             (X10 <= 106)?
               (X3 <= 39)?
                 (X3 <= 18)?
                   (X4 <= 31)?
                    4
                  :
                    8
                :
                  25
              :
                 (X10 <= 61)?
                  2
                :
                  4
            :
               (X5 <= 83)?
                 (X2 <= 18)?
                   (X2 <= 5)?
                    1
                  :
                    2
                :
                  2
              :
                1
          :
             (X7 <= 152)?
               (X0 <= 85)?
                 (X1 <= 50)?
                   (X10 <= 65)?
                    1
                  :
                    4
                :
                   (X2 <= 17)?
                     (X5 <= 121)?
                       (X0 <= 75)?
                        19
                      :
                        1
                    :
                      2
                  :
                     (X2 <= 59)?
                       (X9 <= 41)?
                        8
                      :
                         (X6 <= 31)?
                          1
                        :
                          2
                    :
                       (X9 <= 44)?
                         (X5 <= 52)?
                           (X3 <= 25)?
                            4
                          :
                            3
                        :
                          9
                      :
                        2
              :
                 (X0 <= 89)?
                  1
                :
                  6
            :
              10
      :
         (X1 <= 78)?
           (X3 <= 68)?
             (X2 <= 172)?
               (X0 <= 6)?
                1
              :
                 (X4 <= 5)?
                  2
                :
                   (X6 <= 21)?
                     (X0 <= 101)?
                       (X0 <= 89)?
                         (X6 <= 2)?
                          1
                        :
                           (X6 <= 20)?
                            9
                          :
                             (X7 <= 66)?
                              1
                            :
                              1
                      :
                        3
                    :
                      8
                  :
                    20
            :
               (X8 <= 93)?
                1
              :
                1
          :
             (X2 <= 104)?
               (X7 <= 101)?
                1
              :
                2
            :
              5
        :
           (X7 <= 70)?
             (X8 <= 213)?
               (X2 <= 12)?
                 (X9 <= 28)?
                  3
                :
                  2
              :
                6
            :
              2
          :
             (X1 <= 116)?
               (X1 <= 84)?
                1
              :
                 (X4 <= 21)?
                  1
                :
                  7
            :
               (X1 <= 123)?
                1
              :
                1
    :
       (X10 <= 120)?
         (X1 <= 51)?
           (X6 <= 47)?
             (X8 <= 104)?
               (X0 <= 67)?
                 (X7 <= 87)?
                   (X10 <= 116)?
                    1
                  :
                    1
                :
                  2
              :
                 (X2 <= 165)?
                   (X3 <= 35)?
                     (X3 <= 29)?
                       (X6 <= 13)?
                         (X10 <= 85)?
                          7
                        :
                           (X1 <= 27)?
                            1
                          :
                            3
                      :
                         (X0 <= 100)?
                          3
                        :
                           (X7 <= 163)?
                             (X7 <= 118)?
                               (X2 <= 116)?
                                3
                              :
                                2
                            :
                              11
                          :
                            1
                    :
                       (X8 <= 73)?
                        1
                      :
                        1
                  :
                    6
                :
                  5
            :
               (X5 <= 34)?
                 (X9 <= 71)?
                   (X2 <= 95)?
                    3
                  :
                     (X2 <= 118)?
                       (X6 <= 5)?
                        1
                      :
                         (X6 <= 15)?
                           (X4 <= 33)?
                            2
                          :
                            1
                        :
                          2
                    :
                      5
                :
                   (X2 <= 140)?
                    8
                  :
                    1
              :
                 (X9 <= 62)?
                  10
                :
                   (X7 <= 106)?
                    5
                  :
                     (X7 <= 156)?
                       (X1 <= 28)?
                         (X10 <= 81)?
                          2
                        :
                          2
                      :
                        6
                    :
                      2
          :
             (X5 <= 121)?
               (X2 <= 143)?
                 (X8 <= 123)?
                  8
                :
                   (X2 <= 118)?
                    5
                  :
                    2
              :
                3
            :
               (X0 <= 82)?
                4
              :
                5
        :
           (X6 <= 63)?
             (X4 <= 35)?
               (X1 <= 91)?
                 (X1 <= 63)?
                   (X7 <= 130)?
                     (X7 <= 117)?
                       (X9 <= 71)?
                        8
                      :
                         (X7 <= 96)?
                          2
                        :
                          1
                    :
                      2
                  :
                     (X9 <= 48)?
                      1
                    :
                      12
                :
                   (X0 <= 53)?
                     (X8 <= 182)?
                      17
                    :
                      1
                  :
                     (X1 <= 64)?
                      3
                    :
                       (X8 <= 69)?
                        3
                      :
                         (X8 <= 120)?
                          20
                        :
                           (X2 <= 19)?
                            6
                          :
                            6
              :
                 (X1 <= 93)?
                  4
                :
                   (X10 <= 77)?
                     (X7 <= 142)?
                      5
                    :
                      3
                  :
                     (X1 <= 138)?
                      11
                    :
                      1
            :
               (X6 <= 50)?
                 (X2 <= 59)?
                   (X3 <= 27)?
                    2
                  :
                     (X3 <= 51)?
                       (X3 <= 34)?
                        4
                      :
                         (X5 <= 92)?
                          1
                        :
                          1
                    :
                      1
                :
                   (X2 <= 155)?
                     (X4 <= 55)?
                      12
                    :
                      1
                  :
                    2
              :
                6
          :
             (X9 <= 130)?
               (X2 <= 58)?
                 (X3 <= 22)?
                  1
                :
                   (X10 <= 110)?
                    1
                  :
                    1
              :
                15
            :
              4
      :
         (X10 <= 179)?
           (X9 <= 56)?
             (X6 <= 9)?
               (X3 <= 18)?
                1
              :
                6
            :
               (X3 <= 20)?
                 (X2 <= 104)?
                  1
                :
                  1
              :
                 (X0 <= 177)?
                   (X9 <= 54)?
                    14
                  :
                    1
                :
                  1
          :
             (X5 <= 49)?
               (X9 <= 79)?
                 (X0 <= 127)?
                  22
                :
                   (X3 <= 29)?
                    1
                  :
                    3
              :
                 (X5 <= 29)?
                   (X1 <= 39)?
                    1
                  :
                    5
                :
                  3
            :
               (X3 <= 39)?
                 (X10 <= 124)?
                  4
                :
                   (X2 <= 12)?
                    3
                  :
                     (X6 <= 28)?
                      4
                    :
                       (X6 <= 34)?
                        3
                      :
                         (X4 <= 18)?
                          2
                        :
                           (X8 <= 120)?
                             (X10 <= 138)?
                              2
                            :
                               (X4 <= 26)?
                                2
                              :
                                1
                          :
                            6
              :
                 (X10 <= 169)?
                  3
                :
                  1
        :
           (X6 <= 44)?
             (X4 <= 19)?
              2
            :
               (X9 <= 67)?
                3
              :
                2
          :
             (X5 <= 83)?
              2
            :
              3
;
endmodule
