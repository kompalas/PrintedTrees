module top(X0, X1, X2, X3, X6, X7, X8, X9, X10, X11, X12, X13, X14, X15, X16, X17, X18, X19, out);
input [7:0] X0;
input [7:0] X1;
input [7:0] X2;
input [7:0] X3;
input [7:0] X6;
input [7:0] X7;
input [7:0] X8;
input [7:0] X9;
input [7:0] X10;
input [7:0] X11;
input [7:0] X12;
input [7:0] X13;
input [7:0] X14;
input [7:0] X15;
input [7:0] X16;
input [7:0] X17;
input [7:0] X18;
input [7:0] X19;
output [1:0] out;
assign out = 
   (X7 <= 162)?
     (X17 <= 86)?
       (X12 <= 47)?
         (X8 <= 222)?
          15
        :
          1
      :
         (X13 <= 57)?
          1
        :
          3
    :
       (X0 <= 149)?
         (X6 <= 26)?
           (X16 <= 86)?
            1
          :
             (X8 <= 24)?
               (X16 <= 160)?
                87
              :
                 (X0 <= 133)?
                   (X1 <= 40)?
                     (X17 <= 150)?
                      1
                    :
                      4
                  :
                    4
                :
                  32
            :
              535
        :
           (X2 <= 9)?
             (X10 <= 65)?
              31
            :
               (X14 <= 28)?
                1
              :
                1
          :
             (X1 <= 34)?
               (X13 <= 105)?
                1
              :
                3
            :
               (X19 <= 57)?
                6
              :
                 (X1 <= 67)?
                  2
                :
                  1
      :
         (X1 <= 20)?
           (X18 <= 173)?
             (X6 <= 26)?
               (X9 <= 165)?
                 (X2 <= 5)?
                  60
                :
                   (X2 <= 20)?
                    2
                  :
                    1
              :
                2
            :
              4
          :
             (X0 <= 187)?
               (X3 <= 111)?
                 (X18 <= 191)?
                  14
                :
                   (X11 <= 46)?
                    2
                  :
                    2
              :
                3
            :
               (X9 <= 172)?
                 (X13 <= 98)?
                   (X3 <= 43)?
                     (X15 <= 13)?
                      3
                    :
                       (X16 <= 199)?
                        1
                      :
                        1
                  :
                    16
                :
                   (X0 <= 232)?
                     (X7 <= 121)?
                       (X12 <= 189)?
                        4
                      :
                         (X1 <= 7)?
                          3
                        :
                          1
                    :
                      6
                  :
                     (X1 <= 7)?
                      6
                    :
                      1
              :
                4
        :
           (X3 <= 43)?
             (X9 <= 27)?
               (X19 <= 1)?
                2
              :
                33
            :
               (X10 <= 23)?
                1
              :
                3
          :
             (X15 <= 38)?
              144
            :
               (X12 <= 178)?
                5
              :
                1
  :
     (X9 <= 18)?
       (X17 <= 76)?
         (X13 <= 247)?
           (X14 <= 156)?
            45
          :
             (X6 <= 26)?
              1
            :
              1
        :
          2
      :
         (X7 <= 213)?
           (X19 <= 2)?
             (X12 <= 88)?
              5
            :
               (X3 <= 43)?
                 (X7 <= 183)?
                  2
                :
                  4
              :
                22
          :
             (X6 <= 77)?
              112
            :
               (X2 <= 1)?
                3
              :
                2
        :
           (X18 <= 147)?
            5
          :
            3
    :
       (X9 <= 193)?
         (X7 <= 230)?
           (X0 <= 145)?
             (X8 <= 13)?
               (X3 <= 94)?
                 (X1 <= 34)?
                   (X7 <= 227)?
                    26
                  :
                     (X9 <= 117)?
                      1
                    :
                      1
                :
                  2
              :
                 (X14 <= 114)?
                  4
                :
                  1
            :
               (X14 <= 78)?
                16
              :
                2
          :
             (X9 <= 77)?
               (X7 <= 193)?
                 (X9 <= 75)?
                   (X16 <= 210)?
                    37
                  :
                     (X1 <= 7)?
                      2
                    :
                      1
                :
                  1
              :
                 (X13 <= 93)?
                   (X2 <= 1)?
                    4
                  :
                    3
                :
                  4
            :
              82
        :
           (X3 <= 51)?
            8
          :
            2
      :
         (X3 <= 85)?
          24
        :
           (X8 <= 9)?
            1
          :
            2
;
endmodule
