module top(X0, X1, X2, X3, out);
input [7:0] X0;
input [7:0] X1;
input [7:0] X2;
input [7:0] X3;
output [1:0] out;
assign out = 
   (X0[7:6] <= 0)?
     (X2[7:6] <= 0)?
       (X1[7:5] <= 0)?
         (X3[7:6] <= 0)?
          2
        :
           (X0[7:6] <= 0)?
            4
          :
             (X3[7:6] <= 0)?
               (X1[7:5] <= 0)?
                 (X3[7:6] <= 0)?
                  1
                :
                  1
              :
                2
            :
               (X3[7:6] <= 1)?
                 (X1[7:4] <= 0)?
                  1
                :
                  1
              :
                2
      :
         (X3[7:5] <= 5)?
           (X3[7:6] <= 0)?
            11
          :
             (X0[7:5] <= 0)?
               (X1[7:4] <= 13)?
                1
              :
                1
            :
              3
        :
           (X1[7:6] <= 1)?
            1
          :
            2
    :
       (X3[7:6] <= 0)?
         (X1[7:6] <= 1)?
           (X2[7:6] <= 0)?
             (X0[7:6] <= 0)?
               (X3[7:5] <= 0)?
                 (X1[7:6] <= 0)?
                  1
                :
                  2
              :
                5
            :
               (X1[7:6] <= 0)?
                2
              :
                 (X3[7:6] <= 0)?
                  3
                :
                   (X2[7:6] <= 0)?
                     (X1[7:6] <= 0)?
                      1
                    :
                      1
                  :
                     (X1[7:6] <= 2)?
                      1
                    :
                      1
          :
             (X3[7:4] <= 0)?
               (X0[7:6] <= 0)?
                4
              :
                 (X2[7:6] <= 0)?
                  1
                :
                  2
            :
              11
        :
           (X2[7:5] <= 5)?
             (X0[7:6] <= 0)?
               (X3[7:6] <= 0)?
                3
              :
                1
            :
              5
          :
             (X3[7:6] <= 0)?
               (X0[7:5] <= 0)?
                 (X1[7:5] <= 7)?
                   (X2[7:6] <= 3)?
                    1
                  :
                    1
                :
                   (X2[7:6] <= 0)?
                    1
                  :
                    1
              :
                3
            :
               (X0[7:6] <= 0)?
                4
              :
                 (X2[7:6] <= 1)?
                  1
                :
                   (X1[7:6] <= 1)?
                    1
                  :
                    1
      :
         (X1[7:6] <= 1)?
          72
        :
           (X2[7:4] <= 3)?
             (X0[7:6] <= 0)?
              2
            :
               (X3[7:6] <= 1)?
                1
              :
                1
          :
            10
  :
     (X3[7:6] <= 1)?
       (X1[7:6] <= 0)?
         (X2[7:6] <= 0)?
           (X0[7:6] <= 0)?
             (X2[7:6] <= 0)?
              1
            :
              1
          :
            6
        :
           (X3[7:6] <= 0)?
             (X0[7:6] <= 1)?
              1
            :
               (X2[7:4] <= 7)?
                2
              :
                 (X2[7:4] <= 10)?
                   (X0[7:6] <= 0)?
                    1
                  :
                    1
                :
                  1
          :
            8
      :
         (X2[7:6] <= 0)?
          46
        :
           (X3[7:6] <= 0)?
            20
          :
             (X1[7:6] <= 0)?
               (X0[7:6] <= 4)?
                 (X2[7:6] <= 2)?
                   (X0[7:5] <= 4)?
                    1
                  :
                    1
                :
                  1
              :
                1
            :
               (X0[7:6] <= 0)?
                 (X2[7:6] <= 1)?
                  3
                :
                  1
              :
                10
    :
       (X2[7:6] <= 0)?
         (X1[7:6] <= 1)?
           (X2[7:6] <= 0)?
             (X1[7:6] <= 0)?
               (X0[7:6] <= 2)?
                2
              :
                 (X3[7:6] <= 0)?
                  2
                :
                   (X0[7:6] <= 1)?
                    1
                  :
                     (X3[7:6] <= 1)?
                      1
                    :
                      1
            :
              7
          :
             (X1[7:5] <= 0)?
              6
            :
               (X3[7:6] <= 3)?
                 (X0[7:6] <= 0)?
                  1
                :
                   (X0[7:6] <= 1)?
                     (X3[7:6] <= 0)?
                      1
                    :
                      1
                  :
                    1
              :
                 (X0[7:6] <= 3)?
                  2
                :
                  1
        :
           (X0[7:6] <= 0)?
             (X3[7:6] <= 1)?
              7
            :
               (X2[7:6] <= 0)?
                2
              :
                1
          :
            25
      :
         (X1[7:4] <= 5)?
           (X0[7:5] <= 3)?
             (X1[7:6] <= 0)?
              28
            :
               (X3[7:6] <= 0)?
                 (X2[7:6] <= 4)?
                  2
                :
                  2
              :
                7
          :
             (X2[7:6] <= 0)?
               (X3[7:6] <= 0)?
                1
              :
                 (X1[7:6] <= 1)?
                  2
                :
                  1
            :
              13
        :
           (X2[7:6] <= 0)?
             (X0[7:6] <= 0)?
               (X3[7:6] <= 0)?
                3
              :
                1
            :
              7
          :
             (X3[7:5] <= 3)?
               (X0[7:6] <= 4)?
                 (X1[7:5] <= 3)?
                   (X2[7:6] <= 2)?
                    1
                  :
                    1
                :
                  1
              :
                6
            :
               (X0[7:4] <= 7)?
                6
              :
                 (X2[7:6] <= 2)?
                   (X1[7:6] <= 1)?
                     (X3[7:6] <= 4)?
                       (X0[7:6] <= 3)?
                        1
                      :
                        1
                    :
                       (X0[7:5] <= 3)?
                        1
                      :
                        1
                  :
                    2
                :
                   (X3[7:6] <= 2)?
                     (X0[7:6] <= 2)?
                      1
                    :
                      1
                  :
                    2
;
endmodule
