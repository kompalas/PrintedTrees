module top(X0, X1, X6, X9, X12, X13, X18, X20, X23, X28, X30, X32, X36, X37, X38, X40, X42, X49, X50, X51, X52, X53, X54, X55, X56, X57, X59, X62, X63, X65, X69, X71, X73, X76, X78, X86, X89, X98, X99, X100, X101, X102, X106, X110, X118, X120, X121, X133, X135, X138, X139, X140, X142, X147, X149, X156, X158, X159, X161, X166, X167, X168, X177, X181, X183, X184, X186, X187, X188, X190, X194, X197, X198, X199, X207, X211, X228, X230, X237, X239, X242, X249, X263, X271, X276, X289, X291, X292, X301, X304, X305, X309, X317, X322, X323, X327, X330, X331, X334, X335, X354, X361, X363, X368, X371, X373, X377, X381, X382, X384, X394, X397, X410, X412, X423, X427, X429, X435, X446, X451, X452, X455, X457, X460, X472, X479, X481, X488, X493, X497, X505, X509, X514, X522, X538, X551, X553, X554, X558, X559, X560, out);
input [7:0] X0;
input [7:0] X1;
input [7:0] X6;
input [7:0] X9;
input [7:0] X12;
input [7:0] X13;
input [7:0] X18;
input [7:0] X20;
input [7:0] X23;
input [7:0] X28;
input [7:0] X30;
input [7:0] X32;
input [7:0] X36;
input [7:0] X37;
input [7:0] X38;
input [7:0] X40;
input [7:0] X42;
input [7:0] X49;
input [7:0] X50;
input [7:0] X51;
input [7:0] X52;
input [7:0] X53;
input [7:0] X54;
input [7:0] X55;
input [7:0] X56;
input [7:0] X57;
input [7:0] X59;
input [7:0] X62;
input [7:0] X63;
input [7:0] X65;
input [7:0] X69;
input [7:0] X71;
input [7:0] X73;
input [7:0] X76;
input [7:0] X78;
input [7:0] X86;
input [7:0] X89;
input [7:0] X98;
input [7:0] X99;
input [7:0] X100;
input [7:0] X101;
input [7:0] X102;
input [7:0] X106;
input [7:0] X110;
input [7:0] X118;
input [7:0] X120;
input [7:0] X121;
input [7:0] X133;
input [7:0] X135;
input [7:0] X138;
input [7:0] X139;
input [7:0] X140;
input [7:0] X142;
input [7:0] X147;
input [7:0] X149;
input [7:0] X156;
input [7:0] X158;
input [7:0] X159;
input [7:0] X161;
input [7:0] X166;
input [7:0] X167;
input [7:0] X168;
input [7:0] X177;
input [7:0] X181;
input [7:0] X183;
input [7:0] X184;
input [7:0] X186;
input [7:0] X187;
input [7:0] X188;
input [7:0] X190;
input [7:0] X194;
input [7:0] X197;
input [7:0] X198;
input [7:0] X199;
input [7:0] X207;
input [7:0] X211;
input [7:0] X228;
input [7:0] X230;
input [7:0] X237;
input [7:0] X239;
input [7:0] X242;
input [7:0] X249;
input [7:0] X263;
input [7:0] X271;
input [7:0] X276;
input [7:0] X289;
input [7:0] X291;
input [7:0] X292;
input [7:0] X301;
input [7:0] X304;
input [7:0] X305;
input [7:0] X309;
input [7:0] X317;
input [7:0] X322;
input [7:0] X323;
input [7:0] X327;
input [7:0] X330;
input [7:0] X331;
input [7:0] X334;
input [7:0] X335;
input [7:0] X354;
input [7:0] X361;
input [7:0] X363;
input [7:0] X368;
input [7:0] X371;
input [7:0] X373;
input [7:0] X377;
input [7:0] X381;
input [7:0] X382;
input [7:0] X384;
input [7:0] X394;
input [7:0] X397;
input [7:0] X410;
input [7:0] X412;
input [7:0] X423;
input [7:0] X427;
input [7:0] X429;
input [7:0] X435;
input [7:0] X446;
input [7:0] X451;
input [7:0] X452;
input [7:0] X455;
input [7:0] X457;
input [7:0] X460;
input [7:0] X472;
input [7:0] X479;
input [7:0] X481;
input [7:0] X488;
input [7:0] X493;
input [7:0] X497;
input [7:0] X505;
input [7:0] X509;
input [7:0] X514;
input [7:0] X522;
input [7:0] X538;
input [7:0] X551;
input [7:0] X553;
input [7:0] X554;
input [7:0] X558;
input [7:0] X559;
input [7:0] X560;
output [2:0] out;
assign out = 
   (X102 <= 157)?
     (X56 <= 70)?
       (X63 <= 61)?
         (X133 <= 248)?
           (X242 <= 6)?
            3
          :
             (X121 <= 128)?
              38
            :
              2
        :
          308
      :
         (X54 <= 227)?
           (X42 <= 198)?
             (X133 <= 221)?
              1
            :
              18
          :
             (X98 <= 1)?
              2
            :
              22
        :
           (X139 <= 3)?
             (X363 <= 10)?
              6
            :
              1
          :
            24
    :
       (X460 <= 0)?
         (X40 <= 234)?
          152
        :
           (X289 <= 25)?
             (X55 <= 134)?
               (X460 <= 0)?
                55
              :
                 (X335 <= 0)?
                   (X49 <= 234)?
                     (X42 <= 131)?
                      13
                    :
                      1
                  :
                     (X156 <= 118)?
                       (X188 <= 113)?
                        1
                      :
                        5
                    :
                      14
                :
                  17
            :
               (X559 <= 157)?
                 (X410 <= 0)?
                  41
                :
                   (X488 <= 0)?
                    3
                  :
                    1
              :
                6
          :
             (X110 <= 99)?
               (X78 <= 199)?
                5
              :
                2
            :
              75
      :
         (X51 <= 104)?
           (X239 <= 56)?
             (X50 <= 138)?
               (X49 <= 216)?
                8
              :
                 (X49 <= 238)?
                   (X554 <= 112)?
                     (X30 <= 125)?
                       (X138 <= 0)?
                        1
                      :
                        2
                    :
                      16
                  :
                    262
                :
                   (X455 <= 40)?
                     (X57 <= 3)?
                       (X159 <= 182)?
                        11
                      :
                        2
                    :
                       (X554 <= 186)?
                        10
                      :
                        1
                  :
                    32
            :
               (X57 <= 13)?
                 (X168 <= 10)?
                   (X106 <= 162)?
                     (X323 <= 1)?
                      1
                    :
                      3
                  :
                    24
                :
                  5
              :
                 (X435 <= 15)?
                  42
                :
                  2
          :
             (X76 <= 241)?
              3
            :
               (X140 <= 72)?
                1
              :
                1
        :
           (X57 <= 12)?
             (X230 <= 17)?
               (X32 <= 132)?
                 (X331 <= 0)?
                   (X52 <= 254)?
                     (X184 <= 112)?
                      60
                    :
                      2
                  :
                    4
                :
                   (X228 <= 8)?
                    10
                  :
                     (X497 <= 0)?
                      16
                    :
                       (X481 <= 1)?
                        6
                      :
                        2
              :
                 (X69 <= 49)?
                   (X147 <= 99)?
                     (X301 <= 157)?
                      7
                    :
                      1
                  :
                     (X309 <= 1)?
                      24
                    :
                       (X161 <= 87)?
                        3
                      :
                        3
                :
                   (X371 <= 133)?
                     (X36 <= 92)?
                       (X551 <= 166)?
                        3
                      :
                        1
                    :
                       (X194 <= 99)?
                         (X101 <= 3)?
                          2
                        :
                          2
                      :
                        53
                  :
                     (X40 <= 247)?
                       (X158 <= 197)?
                        9
                      :
                        1
                    :
                      7
            :
               (X457 <= 62)?
                3
              :
                 (X86 <= 37)?
                  1
                :
                  2
          :
             (X446 <= 163)?
              59
            :
              2
  :
     (X65 <= 81)?
       (X69 <= 62)?
         (X560 <= 132)?
           (X371 <= 91)?
             (X335 <= 26)?
              2
            :
              5
          :
             (X493 <= 48)?
              7
            :
               (X384 <= 7)?
                1
              :
                2
        :
           (X330 <= 6)?
             (X71 <= 36)?
              4
            :
               (X429 <= 72)?
                19
              :
                1
          :
             (X381 <= 5)?
               (X20 <= 49)?
                7
              :
                 (X142 <= 152)?
                  2
                :
                  1
            :
               (X412 <= 16)?
                 (X6 <= 35)?
                  4
                :
                   (X199 <= 80)?
                     (X317 <= 18)?
                      9
                    :
                      4
                  :
                     (X382 <= 6)?
                      1
                    :
                      144
              :
                 (X559 <= 99)?
                  8
                :
                   (X451 <= 93)?
                     (X354 <= 69)?
                      4
                    :
                       (X228 <= 102)?
                        2
                      :
                        1
                  :
                     (X40 <= 244)?
                      24
                    :
                      3
      :
         (X330 <= 10)?
           (X42 <= 68)?
            6
          :
             (X135 <= 88)?
               (X166 <= 127)?
                 (X0 <= 139)?
                  2
                :
                   (X373 <= 24)?
                    1
                  :
                    133
              :
                2
            :
               (X553 <= 47)?
                14
              :
                8
        :
           (X89 <= 90)?
             (X57 <= 3)?
               (X538 <= 157)?
                 (X158 <= 174)?
                   (X304 <= 11)?
                    2
                  :
                    12
                :
                   (X479 <= 2)?
                    3
                  :
                    7
              :
                20
            :
               (X38 <= 115)?
                 (X37 <= 207)?
                   (X472 <= 40)?
                     (X505 <= 22)?
                       (X211 <= 144)?
                        4
                      :
                        4
                    :
                       (X237 <= 172)?
                        88
                      :
                        1
                  :
                     (X149 <= 84)?
                      6
                    :
                       (X99 <= 103)?
                        6
                      :
                        2
                :
                   (X177 <= 13)?
                    5
                  :
                    1
              :
                 (X167 <= 64)?
                   (X368 <= 154)?
                    3
                  :
                    22
                :
                   (X18 <= 14)?
                    4
                  :
                    5
          :
             (X427 <= 63)?
               (X514 <= 114)?
                65
              :
                 (X249 <= 135)?
                  5
                :
                  3
            :
               (X558 <= 20)?
                 (X292 <= 12)?
                  3
                :
                  11
              :
                 (X73 <= 55)?
                   (X186 <= 149)?
                    12
                  :
                    1
                :
                   (X23 <= 118)?
                     (X334 <= 30)?
                      1
                    :
                      4
                  :
                    16
    :
       (X509 <= 79)?
         (X55 <= 179)?
           (X42 <= 131)?
             (X100 <= 102)?
               (X305 <= 43)?
                 (X460 <= 4)?
                   (X28 <= 121)?
                     (X190 <= 133)?
                      1
                    :
                      1
                  :
                    11
                :
                   (X452 <= 83)?
                     (X538 <= 85)?
                      5
                    :
                       (X50 <= 123)?
                        11
                      :
                        3
                  :
                     (X197 <= 119)?
                       (X52 <= 246)?
                         (X12 <= 172)?
                           (X271 <= 91)?
                            9
                          :
                            2
                        :
                           (X59 <= 1)?
                            2
                          :
                            8
                      :
                         (X242 <= 53)?
                           (X522 <= 78)?
                             (X207 <= 13)?
                              1
                            :
                              6
                          :
                            10
                        :
                          23
                    :
                       (X23 <= 184)?
                         (X228 <= 108)?
                           (X263 <= 133)?
                            123
                          :
                             (X291 <= 18)?
                              2
                            :
                              5
                        :
                           (X423 <= 77)?
                            5
                          :
                             (X377 <= 125)?
                              15
                            :
                              1
                      :
                        4
              :
                 (X322 <= 21)?
                  18
                :
                   (X13 <= 156)?
                    1
                  :
                    2
            :
               (X371 <= 71)?
                 (X118 <= 116)?
                   (X361 <= 80)?
                    2
                  :
                    2
                :
                  5
              :
                 (X1 <= 141)?
                  144
                :
                   (X551 <= 138)?
                    2
                  :
                    6
          :
             (X49 <= 228)?
               (X69 <= 43)?
                1
              :
                5
            :
              14
        :
           (X53 <= 154)?
             (X181 <= 76)?
               (X89 <= 52)?
                 (X327 <= 5)?
                  2
                :
                  3
              :
                52
            :
               (X198 <= 178)?
                 (X394 <= 46)?
                  9
                :
                  1
              :
                23
          :
             (X488 <= 4)?
               (X187 <= 170)?
                9
              :
                 (X120 <= 112)?
                  1
                :
                  1
            :
              34
      :
         (X57 <= 9)?
           (X55 <= 171)?
             (X9 <= 80)?
              3
            :
              72
          :
            5
        :
           (X276 <= 50)?
             (X53 <= 75)?
              5
            :
               (X183 <= 200)?
                 (X397 <= 38)?
                   (X317 <= 25)?
                    1
                  :
                    1
                :
                  2
              :
                24
          :
             (X62 <= 65)?
              2
            :
              13
;
endmodule
