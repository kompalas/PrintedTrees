module top(X16, out);
input [7:0] X16;
output [3:0] out;
assign out = 
   (X16[7:5] <= 0)?
    800
  :
     (X16[7:1] <= 19)?
      794
    :
       (X16[7:6] <= 1)?
        793
      :
         (X16[7:3] <= 23)?
           (X16[7:2] <= 31)?
             (X16[7:4] <= 7)?
              734
            :
              786
          :
             (X16[7:5] <= 6)?
              738
            :
              752
        :
           (X16 <= 212)?
            805
          :
             (X16[7:2] <= 61)?
              747
            :
              745
;
endmodule
