module top(X0, X1, X6, X9, X12, X13, X18, X20, X23, X28, X30, X32, X36, X37, X38, X40, X42, X49, X50, X51, X52, X53, X54, X55, X56, X57, X59, X62, X63, X65, X69, X71, X73, X76, X78, X86, X89, X98, X99, X100, X101, X102, X106, X110, X118, X120, X121, X133, X135, X138, X139, X140, X142, X147, X149, X156, X158, X159, X161, X166, X167, X168, X177, X181, X183, X184, X186, X187, X188, X190, X194, X197, X198, X199, X207, X211, X228, X230, X237, X239, X242, X249, X263, X271, X276, X289, X291, X292, X301, X304, X305, X309, X317, X322, X323, X327, X330, X331, X334, X335, X354, X361, X363, X368, X371, X373, X377, X381, X382, X384, X394, X397, X410, X412, X423, X427, X429, X435, X446, X451, X452, X455, X457, X460, X472, X479, X481, X488, X493, X497, X505, X509, X514, X522, X538, X551, X553, X554, X558, X559, X560, out);
input [7:0] X0;
input [7:0] X1;
input [7:0] X6;
input [7:0] X9;
input [7:0] X12;
input [7:0] X13;
input [7:0] X18;
input [7:0] X20;
input [7:0] X23;
input [7:0] X28;
input [7:0] X30;
input [7:0] X32;
input [7:0] X36;
input [7:0] X37;
input [7:0] X38;
input [7:0] X40;
input [7:0] X42;
input [7:0] X49;
input [7:0] X50;
input [7:0] X51;
input [7:0] X52;
input [7:0] X53;
input [7:0] X54;
input [7:0] X55;
input [7:0] X56;
input [7:0] X57;
input [7:0] X59;
input [7:0] X62;
input [7:0] X63;
input [7:0] X65;
input [7:0] X69;
input [7:0] X71;
input [7:0] X73;
input [7:0] X76;
input [7:0] X78;
input [7:0] X86;
input [7:0] X89;
input [7:0] X98;
input [7:0] X99;
input [7:0] X100;
input [7:0] X101;
input [7:0] X102;
input [7:0] X106;
input [7:0] X110;
input [7:0] X118;
input [7:0] X120;
input [7:0] X121;
input [7:0] X133;
input [7:0] X135;
input [7:0] X138;
input [7:0] X139;
input [7:0] X140;
input [7:0] X142;
input [7:0] X147;
input [7:0] X149;
input [7:0] X156;
input [7:0] X158;
input [7:0] X159;
input [7:0] X161;
input [7:0] X166;
input [7:0] X167;
input [7:0] X168;
input [7:0] X177;
input [7:0] X181;
input [7:0] X183;
input [7:0] X184;
input [7:0] X186;
input [7:0] X187;
input [7:0] X188;
input [7:0] X190;
input [7:0] X194;
input [7:0] X197;
input [7:0] X198;
input [7:0] X199;
input [7:0] X207;
input [7:0] X211;
input [7:0] X228;
input [7:0] X230;
input [7:0] X237;
input [7:0] X239;
input [7:0] X242;
input [7:0] X249;
input [7:0] X263;
input [7:0] X271;
input [7:0] X276;
input [7:0] X289;
input [7:0] X291;
input [7:0] X292;
input [7:0] X301;
input [7:0] X304;
input [7:0] X305;
input [7:0] X309;
input [7:0] X317;
input [7:0] X322;
input [7:0] X323;
input [7:0] X327;
input [7:0] X330;
input [7:0] X331;
input [7:0] X334;
input [7:0] X335;
input [7:0] X354;
input [7:0] X361;
input [7:0] X363;
input [7:0] X368;
input [7:0] X371;
input [7:0] X373;
input [7:0] X377;
input [7:0] X381;
input [7:0] X382;
input [7:0] X384;
input [7:0] X394;
input [7:0] X397;
input [7:0] X410;
input [7:0] X412;
input [7:0] X423;
input [7:0] X427;
input [7:0] X429;
input [7:0] X435;
input [7:0] X446;
input [7:0] X451;
input [7:0] X452;
input [7:0] X455;
input [7:0] X457;
input [7:0] X460;
input [7:0] X472;
input [7:0] X479;
input [7:0] X481;
input [7:0] X488;
input [7:0] X493;
input [7:0] X497;
input [7:0] X505;
input [7:0] X509;
input [7:0] X514;
input [7:0] X522;
input [7:0] X538;
input [7:0] X551;
input [7:0] X553;
input [7:0] X554;
input [7:0] X558;
input [7:0] X559;
input [7:0] X560;
output [2:0] out;
assign out = 
   (X102[7:3] <= 21)?
     (X56 <= 73)?
       (X63[7:1] <= 35)?
         (X133[7:1] <= 123)?
           (X242[7:5] <= 2)?
            3
          :
             (X121[7:1] <= 66)?
              38
            :
              2
        :
          308
      :
         (X54[7:1] <= 114)?
           (X42[7:1] <= 101)?
             (X133[7:2] <= 57)?
              1
            :
              18
          :
             (X98[7:2] <= 4)?
              2
            :
              22
        :
           (X139[7:1] <= 6)?
             (X363[7:1] <= 8)?
              6
            :
              1
          :
            24
    :
       (X460[7:2] <= 0)?
         (X40[7:1] <= 117)?
          152
        :
           (X289[7:5] <= 3)?
             (X55[7:4] <= 8)?
               (X460[7:1] <= 3)?
                55
              :
                 (X335[7:2] <= 1)?
                   (X49[7:1] <= 118)?
                     (X42[7:2] <= 37)?
                      13
                    :
                      1
                  :
                     (X156[7:5] <= 7)?
                       (X188[7:2] <= 31)?
                        1
                      :
                        5
                    :
                      14
                :
                  17
            :
               (X559[7:3] <= 18)?
                 (X410[7:2] <= 2)?
                  41
                :
                   (X488[7:2] <= 0)?
                    3
                  :
                    1
              :
                6
          :
             (X110[7:5] <= 3)?
               (X78[7:5] <= 8)?
                5
              :
                2
            :
              75
      :
         (X51[7:2] <= 30)?
           (X239[7:2] <= 17)?
             (X50[7:2] <= 36)?
               (X49[7:2] <= 55)?
                8
              :
                 (X49[7:3] <= 32)?
                   (X554[7:2] <= 28)?
                     (X30[7:4] <= 9)?
                       (X138[7:3] <= 3)?
                        1
                      :
                        2
                    :
                      16
                  :
                    262
                :
                   (X455[7:4] <= 2)?
                     (X57[7:2] <= 1)?
                       (X159[7:4] <= 11)?
                        11
                      :
                        2
                    :
                       (X554[7:2] <= 50)?
                        10
                      :
                        1
                  :
                    32
            :
               (X57[7:1] <= 4)?
                 (X168[7:2] <= 6)?
                   (X106[7:4] <= 10)?
                     (X323[7:4] <= 1)?
                      1
                    :
                      3
                  :
                    24
                :
                  5
              :
                 (X435[7:2] <= 5)?
                  42
                :
                  2
          :
             (X76[7:2] <= 61)?
              3
            :
               (X140[7:1] <= 37)?
                1
              :
                1
        :
           (X57[7:3] <= 3)?
             (X230[7:3] <= 6)?
               (X32[7:1] <= 69)?
                 (X331[7:4] <= 3)?
                   (X52[7:1] <= 128)?
                     (X184[7:5] <= 4)?
                      60
                    :
                      2
                  :
                    4
                :
                   (X228[7:3] <= 4)?
                    10
                  :
                     (X497[7:2] <= 4)?
                      16
                    :
                       (X481[7:4] <= 0)?
                        6
                      :
                        2
              :
                 (X69[7:2] <= 15)?
                   (X147[7:5] <= 3)?
                     (X301[7:4] <= 14)?
                      7
                    :
                      1
                  :
                     (X309 <= 1)?
                      24
                    :
                       (X161[7:1] <= 44)?
                        3
                      :
                        3
                :
                   (X371[7:2] <= 32)?
                     (X36[7:6] <= 1)?
                       (X551[7:2] <= 43)?
                        3
                      :
                        1
                    :
                       (X194[7:2] <= 25)?
                         (X101[7:4] <= 3)?
                          2
                        :
                          2
                      :
                        53
                  :
                     (X40[7:3] <= 32)?
                       (X158[7:5] <= 4)?
                        9
                      :
                        1
                    :
                      7
            :
               (X457[7:3] <= 6)?
                3
              :
                 (X86[7:3] <= 7)?
                  1
                :
                  2
          :
             (X446[7:3] <= 21)?
              59
            :
              2
  :
     (X65[7:3] <= 10)?
       (X69[7:3] <= 8)?
         (X560[7:3] <= 19)?
           (X371[7:3] <= 11)?
             (X335[7:1] <= 12)?
              2
            :
              5
          :
             (X493[7:4] <= 7)?
              7
            :
               (X384[7:1] <= 6)?
                1
              :
                2
        :
           (X330[7:1] <= 5)?
             (X71[7:2] <= 8)?
              4
            :
               (X429[7:1] <= 36)?
                19
              :
                1
          :
             (X381[7:3] <= 1)?
               (X20[7:3] <= 6)?
                7
              :
                 (X142[7:1] <= 79)?
                  2
                :
                  1
            :
               (X412[7:2] <= 6)?
                 (X6[7:3] <= 4)?
                  4
                :
                   (X199[7:3] <= 10)?
                     (X317[7:6] <= 1)?
                      9
                    :
                      4
                  :
                     (X382[7:1] <= 2)?
                      1
                    :
                      144
              :
                 (X559[7:4] <= 8)?
                  8
                :
                   (X451[7:2] <= 25)?
                     (X354[7:5] <= 6)?
                      4
                    :
                       (X228[7:4] <= 8)?
                        2
                      :
                        1
                  :
                     (X40[7:5] <= 8)?
                      24
                    :
                      3
      :
         (X330[7:1] <= 6)?
           (X42[7:1] <= 38)?
            6
          :
             (X135[7:4] <= 8)?
               (X166[7:1] <= 67)?
                 (X0[7:3] <= 15)?
                  2
                :
                   (X373[7:1] <= 14)?
                    1
                  :
                    133
              :
                2
            :
               (X553[7:4] <= 6)?
                14
              :
                8
        :
           (X89[7:5] <= 3)?
             (X57[7:1] <= 5)?
               (X538[7:1] <= 79)?
                 (X158[7:2] <= 47)?
                   (X304[7:1] <= 5)?
                    2
                  :
                    12
                :
                   (X479[7:3] <= 0)?
                    3
                  :
                    7
              :
                20
            :
               (X38[7:2] <= 30)?
                 (X37[7:1] <= 102)?
                   (X472[7:6] <= 4)?
                     (X505[7:2] <= 5)?
                       (X211[7:1] <= 71)?
                        4
                      :
                        4
                    :
                       (X237[7:3] <= 19)?
                        88
                      :
                        1
                  :
                     (X149[7:6] <= 0)?
                      6
                    :
                       (X99[7:2] <= 28)?
                        6
                      :
                        2
                :
                   (X177[7:4] <= 3)?
                    5
                  :
                    1
              :
                 (X167[7:5] <= 2)?
                   (X368[7:3] <= 20)?
                    3
                  :
                    22
                :
                   (X18[7:2] <= 3)?
                    4
                  :
                    5
          :
             (X427[7:4] <= 4)?
               (X514[7:3] <= 13)?
                65
              :
                 (X249[7:5] <= 1)?
                  5
                :
                  3
            :
               (X558[7:5] <= 2)?
                 (X292[7:3] <= 3)?
                  3
                :
                  11
              :
                 (X73[7:4] <= 6)?
                   (X186[7:4] <= 11)?
                    12
                  :
                    1
                :
                   (X23[7:2] <= 28)?
                     (X334[7:2] <= 11)?
                      1
                    :
                      4
                  :
                    16
    :
       (X509[7:6] <= 0)?
         (X55[7:1] <= 91)?
           (X42[7:5] <= 4)?
             (X100[7:1] <= 49)?
               (X305[7:4] <= 6)?
                 (X460[7:1] <= 5)?
                   (X28[7:1] <= 61)?
                     (X190[7:2] <= 38)?
                      1
                    :
                      1
                  :
                    11
                :
                   (X452[7:3] <= 11)?
                     (X538[7:4] <= 6)?
                      5
                    :
                       (X50[7:2] <= 35)?
                        11
                      :
                        3
                  :
                     (X197[7:1] <= 61)?
                       (X52[7:4] <= 16)?
                         (X12[7:1] <= 84)?
                           (X271[7:3] <= 14)?
                            9
                          :
                            2
                        :
                           (X59[7:2] <= 0)?
                            2
                          :
                            8
                      :
                         (X242[7:3] <= 8)?
                           (X522[7:2] <= 22)?
                             (X207[7:2] <= 6)?
                              1
                            :
                              6
                          :
                            10
                        :
                          23
                    :
                       (X23[7:4] <= 11)?
                         (X228[7:3] <= 17)?
                           (X263[7:1] <= 68)?
                            123
                          :
                             (X291[7:5] <= 4)?
                              2
                            :
                              5
                        :
                           (X423[7:4] <= 9)?
                            5
                          :
                             (X377[7:1] <= 64)?
                              15
                            :
                              1
                      :
                        4
              :
                 (X322[7:2] <= 8)?
                  18
                :
                   (X13[7:5] <= 8)?
                    1
                  :
                    2
            :
               (X371[7:2] <= 20)?
                 (X118[7:2] <= 33)?
                   (X361[7:2] <= 19)?
                    2
                  :
                    2
                :
                  5
              :
                 (X1[7:5] <= 7)?
                  144
                :
                   (X551[7:3] <= 17)?
                    2
                  :
                    6
          :
             (X49[7:4] <= 16)?
               (X69[7:1] <= 23)?
                1
              :
                5
            :
              14
        :
           (X53[7:1] <= 75)?
             (X181[7:1] <= 42)?
               (X89[7:4] <= 5)?
                 (X327[7:4] <= 1)?
                  2
                :
                  3
              :
                52
            :
               (X198[7:4] <= 14)?
                 (X394[7:1] <= 23)?
                  9
                :
                  1
              :
                23
          :
             (X488[7:1] <= 3)?
               (X187[7:3] <= 23)?
                9
              :
                 (X120[7:3] <= 17)?
                  1
                :
                  1
            :
              34
      :
         (X57[7:4] <= 5)?
           (X55[7:1] <= 84)?
             (X9[7:3] <= 11)?
              3
            :
              72
          :
            5
        :
           (X276[7:2] <= 17)?
             (X53[7:5] <= 0)?
              5
            :
               (X183[7:1] <= 102)?
                 (X397[7:5] <= 0)?
                   (X317[7:3] <= 4)?
                    1
                  :
                    1
                :
                  2
              :
                24
          :
             (X62[7:1] <= 34)?
              2
            :
              13
;
endmodule
