module top(X0, X1, X4, X9, X12, X28, X30, X32, X37, X38, X41, X42, X44, X49, X51, X52, X54, X55, X56, X57, X58, X62, X63, X65, X69, X73, X90, X93, X101, X102, X106, X113, X114, X115, X118, X125, X128, X133, X136, X137, X139, X141, X142, X147, X148, X155, X159, X161, X162, X165, X169, X170, X172, X180, X181, X185, X190, X192, X198, X199, X209, X210, X227, X238, X240, X244, X245, X248, X258, X259, X263, X265, X268, X270, X273, X274, X275, X276, X283, X286, X287, X290, X296, X300, X301, X302, X310, X312, X313, X319, X320, X323, X324, X326, X327, X330, X331, X335, X336, X340, X342, X358, X361, X362, X370, X371, X376, X380, X387, X388, X394, X395, X403, X405, X409, X410, X414, X428, X432, X434, X435, X445, X449, X452, X455, X457, X458, X460, X462, X477, X481, X483, X488, X489, X498, X504, X509, X514, X524, X527, X535, X537, X539, X542, X550, X554, X558, X560, out);
input [7:0] X0;
input [7:0] X1;
input [7:0] X4;
input [7:0] X9;
input [7:0] X12;
input [7:0] X28;
input [7:0] X30;
input [7:0] X32;
input [7:0] X37;
input [7:0] X38;
input [7:0] X41;
input [7:0] X42;
input [7:0] X44;
input [7:0] X49;
input [7:0] X51;
input [7:0] X52;
input [7:0] X54;
input [7:0] X55;
input [7:0] X56;
input [7:0] X57;
input [7:0] X58;
input [7:0] X62;
input [7:0] X63;
input [7:0] X65;
input [7:0] X69;
input [7:0] X73;
input [7:0] X90;
input [7:0] X93;
input [7:0] X101;
input [7:0] X102;
input [7:0] X106;
input [7:0] X113;
input [7:0] X114;
input [7:0] X115;
input [7:0] X118;
input [7:0] X125;
input [7:0] X128;
input [7:0] X133;
input [7:0] X136;
input [7:0] X137;
input [7:0] X139;
input [7:0] X141;
input [7:0] X142;
input [7:0] X147;
input [7:0] X148;
input [7:0] X155;
input [7:0] X159;
input [7:0] X161;
input [7:0] X162;
input [7:0] X165;
input [7:0] X169;
input [7:0] X170;
input [7:0] X172;
input [7:0] X180;
input [7:0] X181;
input [7:0] X185;
input [7:0] X190;
input [7:0] X192;
input [7:0] X198;
input [7:0] X199;
input [7:0] X209;
input [7:0] X210;
input [7:0] X227;
input [7:0] X238;
input [7:0] X240;
input [7:0] X244;
input [7:0] X245;
input [7:0] X248;
input [7:0] X258;
input [7:0] X259;
input [7:0] X263;
input [7:0] X265;
input [7:0] X268;
input [7:0] X270;
input [7:0] X273;
input [7:0] X274;
input [7:0] X275;
input [7:0] X276;
input [7:0] X283;
input [7:0] X286;
input [7:0] X287;
input [7:0] X290;
input [7:0] X296;
input [7:0] X300;
input [7:0] X301;
input [7:0] X302;
input [7:0] X310;
input [7:0] X312;
input [7:0] X313;
input [7:0] X319;
input [7:0] X320;
input [7:0] X323;
input [7:0] X324;
input [7:0] X326;
input [7:0] X327;
input [7:0] X330;
input [7:0] X331;
input [7:0] X335;
input [7:0] X336;
input [7:0] X340;
input [7:0] X342;
input [7:0] X358;
input [7:0] X361;
input [7:0] X362;
input [7:0] X370;
input [7:0] X371;
input [7:0] X376;
input [7:0] X380;
input [7:0] X387;
input [7:0] X388;
input [7:0] X394;
input [7:0] X395;
input [7:0] X403;
input [7:0] X405;
input [7:0] X409;
input [7:0] X410;
input [7:0] X414;
input [7:0] X428;
input [7:0] X432;
input [7:0] X434;
input [7:0] X435;
input [7:0] X445;
input [7:0] X449;
input [7:0] X452;
input [7:0] X455;
input [7:0] X457;
input [7:0] X458;
input [7:0] X460;
input [7:0] X462;
input [7:0] X477;
input [7:0] X481;
input [7:0] X483;
input [7:0] X488;
input [7:0] X489;
input [7:0] X498;
input [7:0] X504;
input [7:0] X509;
input [7:0] X514;
input [7:0] X524;
input [7:0] X527;
input [7:0] X535;
input [7:0] X537;
input [7:0] X539;
input [7:0] X542;
input [7:0] X550;
input [7:0] X554;
input [7:0] X558;
input [7:0] X560;
output [2:0] out;
assign out = 
   (X102[7:6] <= 2)?
     (X56[7:3] <= 7)?
       (X63[7:6] <= 1)?
         (X118[7:6] <= 0)?
           (X137[7:6] <= 0)?
             (X301[7:5] <= 0)?
               (X310[7:5] <= 0)?
                8
              :
                1
            :
              335
          :
            1
        :
           (X327[7:5] <= 0)?
             (X210[7:6] <= 0)?
              3
            :
              1
          :
            5
      :
         (X58[7:5] <= 0)?
           (X51[7:6] <= 0)?
             (X113[7:6] <= 2)?
              17
            :
              1
          :
             (X198[7:5] <= 0)?
              3
            :
              19
        :
           (X560[7:6] <= 0)?
            6
          :
             (X106[7:5] <= 3)?
              1
            :
              22
    :
       (X560[7:5] <= 5)?
         (X49[7:5] <= 6)?
          184
        :
           (X340[7:6] <= 0)?
             (X445[7:5] <= 0)?
              6
            :
               (X199[7:6] <= 2)?
                24
              :
                3
          :
             (X481[7:6] <= 1)?
               (X63[7:6] <= 0)?
                92
              :
                 (X312[7:6] <= 0)?
                  4
                :
                  9
            :
               (X32[7:6] <= 0)?
                 (X326[7:6] <= 1)?
                  2
                :
                  2
              :
                2
      :
         (X139[7:4] <= 0)?
           (X58[7:4] <= 0)?
             (X403[7:5] <= 0)?
               (X57[7:6] <= 0)?
                 (X361[7:6] <= 0)?
                  11
                :
                  1
              :
                 (X259[7:6] <= 0)?
                  10
                :
                  1
            :
               (X320[7:6] <= 0)?
                80
              :
                 (X286[7:5] <= 0)?
                  6
                :
                   (X118[7:6] <= 0)?
                     (X300[7:6] <= 0)?
                      3
                    :
                      3
                  :
                    29
          :
             (X41[7:6] <= 0)?
              6
            :
               (X142[7:5] <= 0)?
                2
              :
                30
        :
           (X51[7:6] <= 0)?
             (X245[7:6] <= 0)?
               (X42[7:6] <= 0)?
                9
              :
                 (X41[7:5] <= 1)?
                   (X460[7:6] <= 0)?
                     (X125[7:6] <= 0)?
                      12
                    :
                       (X394[7:6] <= 0)?
                        10
                      :
                        2
                  :
                     (X65[7:6] <= 0)?
                       (X558[7:5] <= 0)?
                        6
                      :
                         (X263[7:4] <= 7)?
                          36
                        :
                           (X380[7:6] <= 0)?
                            3
                          :
                            1
                    :
                       (X527[7:6] <= 0)?
                        232
                      :
                         (X388[7:6] <= 0)?
                           (X319[7:6] <= 0)?
                            1
                          :
                            33
                        :
                          2
                :
                   (X57[7:6] <= 0)?
                     (X192[7:6] <= 0)?
                      23
                    :
                      4
                  :
                     (X539[7:6] <= 0)?
                      44
                    :
                      3
            :
               (X488[7:6] <= 0)?
                2
              :
                 (X93[7:6] <= 2)?
                  1
                :
                  1
          :
             (X248[7:6] <= 0)?
               (X498[7:6] <= 0)?
                 (X414[7:5] <= 0)?
                  37
                :
                  1
              :
                 (X275[7:6] <= 0)?
                  7
                :
                  4
            :
               (X101[7:5] <= 2)?
                 (X54[7:6] <= 1)?
                   (X290[7:5] <= 0)?
                     (X161[7:6] <= 0)?
                      5
                    :
                       (X190[7:6] <= 2)?
                        14
                      :
                        2
                  :
                    13
                :
                   (X335[7:6] <= 0)?
                    46
                  :
                     (X169[7:6] <= 0)?
                      5
                    :
                      7
              :
                 (X376[7:6] <= 0)?
                  2
                :
                  2
  :
     (X69[7:5] <= 0)?
       (X302[7:6] <= 0)?
         (X38[7:6] <= 0)?
           (X395[7:5] <= 0)?
             (X268[7:5] <= 0)?
              5
            :
              10
          :
             (X30[7:6] <= 0)?
               (X537[7:6] <= 0)?
                2
              :
                1
            :
              7
        :
           (X455[7:6] <= 1)?
            37
          :
            1
      :
         (X52[7:6] <= 2)?
           (X159[7:6] <= 0)?
             (X371[7:4] <= 2)?
              5
            :
               (X358[7:6] <= 0)?
                10
              :
                3
          :
             (X457[7:5] <= 0)?
               (X41[7:6] <= 0)?
                2
              :
                5
            :
               (X136[7:5] <= 0)?
                 (X240[7:6] <= 0)?
                   (X273[7:4] <= 7)?
                    1
                  :
                    1
                :
                  16
              :
                 (X313[7:6] <= 0)?
                  1
                :
                  3
        :
           (X434[7:6] <= 0)?
             (X73[7:6] <= 0)?
               (X449[7:4] <= 0)?
                 (X287[7:5] <= 2)?
                   (X524[7:3] <= 0)?
                    1
                  :
                    23
                :
                  3
              :
                 (X0[7:6] <= 0)?
                  10
                :
                  2
            :
              30
          :
             (X37[7:6] <= 2)?
               (X457[7:6] <= 0)?
                 (X128[7:6] <= 0)?
                   (X462[7:6] <= 0)?
                    7
                  :
                    3
                :
                   (X192[7:6] <= 1)?
                     (X244[7:5] <= 0)?
                      6
                    :
                      3
                  :
                    59
              :
                113
            :
               (X403[7:6] <= 0)?
                1
              :
                9
    :
       (X509[7:4] <= 5)?
         (X37[7:5] <= 1)?
           (X69[7:4] <= 6)?
             (X394[7:6] <= 0)?
               (X265[7:6] <= 1)?
                 (X90[7:5] <= 0)?
                   (X336[7:6] <= 0)?
                    2
                  :
                     (X4[7:4] <= 1)?
                      1
                    :
                      2
                :
                  50
              :
                 (X54[7:6] <= 0)?
                  12
                :
                   (X49[7:6] <= 2)?
                    8
                  :
                    2
            :
               (X57[7:6] <= 0)?
                 (X209[7:6] <= 0)?
                   (X12[7:6] <= 0)?
                    9
                  :
                     (X312[7:4] <= 0)?
                      4
                    :
                       (X62[7:6] <= 0)?
                        16
                      :
                        2
                :
                   (X428[7:6] <= 0)?
                    1
                  :
                    34
              :
                 (X283[7:6] <= 0)?
                   (X483[7:6] <= 0)?
                     (X1[7:5] <= 4)?
                      4
                    :
                       (X324[7:6] <= 0)?
                        31
                      :
                        1
                  :
                     (X504[7:6] <= 1)?
                      12
                    :
                       (X550[7:6] <= 0)?
                        3
                      :
                        1
                :
                   (X342[7:5] <= 0)?
                     (X181[7:6] <= 0)?
                       (X55[7:6] <= 1)?
                         (X435[7:6] <= 0)?
                           (X535[7:6] <= 0)?
                            8
                          :
                            1
                        :
                           (X258[7:6] <= 0)?
                            5
                          :
                            3
                      :
                        19
                    :
                       (X1[7:5] <= 2)?
                        2
                      :
                        12
                  :
                    31
          :
             (X44[7:5] <= 0)?
               (X488[7:6] <= 0)?
                 (X331[7:6] <= 0)?
                  4
                :
                   (X133[7:6] <= 0)?
                    2
                  :
                     (X57[7:5] <= 0)?
                      1
                    :
                      1
              :
                 (X274[7:4] <= 2)?
                   (X162[7:6] <= 0)?
                    189
                  :
                     (X147[7:5] <= 3)?
                       (X185[7:6] <= 1)?
                        22
                      :
                        1
                    :
                      2
                :
                  2
            :
               (X181[7:6] <= 0)?
                 (X452[7:6] <= 0)?
                   (X276[7:6] <= 0)?
                     (X90[7:5] <= 0)?
                      5
                    :
                       (X165[7:6] <= 0)?
                         (X477[7:6] <= 0)?
                          3
                        :
                          1
                      :
                        10
                  :
                     (X405[7:5] <= 0)?
                       (X409[7:6] <= 0)?
                        8
                      :
                        2
                    :
                      9
                :
                   (X28[7:6] <= 0)?
                     (X141[7:5] <= 0)?
                      1
                    :
                      23
                  :
                    2
              :
                 (X180[7:6] <= 0)?
                  44
                :
                  2
        :
           (X409[7:6] <= 0)?
             (X296[7:5] <= 0)?
               (X452[7:6] <= 0)?
                1
              :
                1
            :
              57
          :
             (X159[7:6] <= 0)?
               (X199[7:5] <= 2)?
                 (X238[7:6] <= 1)?
                  21
                :
                   (X410[7:6] <= 0)?
                     (X115[7:5] <= 3)?
                      3
                    :
                      2
                  :
                     (X458[7:6] <= 0)?
                      1
                    :
                      7
              :
                 (X550[7:6] <= 0)?
                  1
                :
                  13
            :
               (X170[7:5] <= 0)?
                 (X387[7:6] <= 0)?
                  2
                :
                  1
              :
                 (X102[7:6] <= 0)?
                  24
                :
                  1
      :
         (X57[7:6] <= 0)?
           (X514[7:6] <= 0)?
             (X9[7:6] <= 2)?
               (X172[7:6] <= 0)?
                 (X227[7:6] <= 0)?
                  16
                :
                  3
              :
                 (X155[7:5] <= 3)?
                  1
                :
                  6
            :
               (X115[7:6] <= 0)?
                 (X114[7:6] <= 0)?
                  1
                :
                  136
              :
                 (X542[7:6] <= 0)?
                  3
                :
                  2
          :
             (X432[7:4] <= 2)?
               (X170[7:5] <= 0)?
                3
              :
                1
            :
               (X458[7:6] <= 0)?
                1
              :
                20
        :
           (X330[7:5] <= 0)?
             (X489[7:5] <= 0)?
              48
            :
              1
          :
             (X38[7:2] <= 15)?
               (X238[7:5] <= 1)?
                 (X199[7:6] <= 0)?
                  32
                :
                  3
              :
                 (X554[7:5] <= 1)?
                  9
                :
                  2
            :
               (X270[7:6] <= 0)?
                 (X434[7:6] <= 0)?
                   (X185[7:6] <= 0)?
                     (X323[7:6] <= 0)?
                      2
                    :
                      8
                  :
                     (X148[7:3] <= 4)?
                      1
                    :
                      6
                :
                   (X370[7:6] <= 0)?
                    12
                  :
                    3
              :
                 (X362[7:6] <= 0)?
                  27
                :
                  1
;
endmodule
