module top(X16, out);
input [7:0] X16;
output [3:0] out;
assign out = 
   (X16 <= 14)?
    796
  :
     (X16 <= 71)?
       (X16 <= 43)?
        785
      :
        815
    :
       (X16 <= 185)?
         (X16 <= 128)?
           (X16 <= 100)?
            711
          :
            799
        :
           (X16 <= 156)?
            749
          :
            752
      :
         (X16 <= 213)?
          831
        :
           (X16 <= 242)?
            747
          :
            709
;
endmodule
