module top(X0, X1, X2, X3, X4, X5, out);
input [7:0] X0;
input [7:0] X1;
input [7:0] X2;
input [7:0] X3;
input [7:0] X4;
input [7:0] X5;
output [1:0] out;
assign out = 
   (X5[7:2] <= 3)?
     (X3[7:5] <= 2)?
       (X4[7:1] <= 66)?
        13
      :
         (X1[7:4] <= 5)?
           (X0[7:2] <= 4)?
            1
          :
            11
        :
           (X4[7:3] <= 21)?
             (X1[7:3] <= 14)?
               (X0[7:4] <= 2)?
                 (X5[7:3] <= 1)?
                  8
                :
                   (X4[7:3] <= 19)?
                    1
                  :
                    1
              :
                 (X3[7:3] <= 6)?
                  3
                :
                   (X0[7:4] <= 3)?
                    1
                  :
                    4
            :
              6
          :
             (X5[7:2] <= 5)?
               (X1[7:3] <= 16)?
                7
              :
                1
            :
              2
    :
       (X4[7:4] <= 8)?
         (X3[7:3] <= 11)?
           (X1[7:2] <= 37)?
             (X4 <= 110)?
              6
            :
               (X5[7:2] <= 2)?
                 (X5[7:4] <= 0)?
                  1
                :
                  3
              :
                3
          :
             (X2 <= 90)?
              1
            :
              2
        :
           (X0[7:4] <= 7)?
             (X0[7:4] <= 7)?
              2
            :
              2
          :
            5
      :
        29
  :
     (X5[7:3] <= 3)?
       (X5[7:2] <= 6)?
         (X4[7:3] <= 23)?
          24
        :
           (X2[7:2] <= 21)?
            3
          :
            1
      :
        1
    :
      75
;
endmodule
